//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "RS_nor.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(144,216)(177,216){1}
reg w1;    //: /sn:0 {0}(140,335)(173,335)(173,384)(216,384){1}
wire w6;    //: /sn:0 {0}(143,426)(158,426)(158,347){1}
//: {2}(160,345)(170,345)(170,389)(216,389){3}
//: {4}(158,343)(158,221)(177,221){5}
wire w4;    //: /sn:0 {0}(198,219)(255,219)(255,216)(286,216){1}
wire w8;    //: /sn:0 {0}(304,382)(276,382)(276,300)(321,300)(321,223){1}
//: {2}(323,221)(442,221)(442,211){3}
//: {4}(319,221)(311,221)(311,219)(307,219){5}
wire w2;    //: /sn:0 {0}(304,387)(237,387){1}
wire w10;    //: /sn:0 {0}(325,385)(357,385){1}
//: {2}(361,385)(443,385)(443,353){3}
//: {4}(359,383)(359,274)(276,274)(276,221)(286,221){5}
//: enddecls

  //: comment g8 @(541,191) /sn:0
  //: /line:"S  R   Q  Q'"
  //: /line:"1  0   1  0"
  //: /line:"0  0   1  0"
  //: /line:"0  1   0  1"
  //: /line:"0  0   0  1"
  //: /line:"1  1   0  0"
  //: /end
  //: joint g4 (w8) @(321, 221) /w:[ 2 -1 4 1 ]
  //: comment g13 @(439,309) /sn:0
  //: /line:"--"
  //: /line:"Q"
  //: /line:""
  //: /end
  _GGAND2 #(6) g2 (.I0(w0), .I1(w6), .Z(w4));   //: @(188,219) /sn:0 /w:[ 1 5 0 ]
  //: SWITCH g1 (w1) @(123,335) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: comment g11 @(228,318) /sn:0
  //: /line:"Set"
  //: /end
  _GGAND2 #(6) g16 (.I0(w1), .I1(w6), .Z(w2));   //: @(227,387) /sn:0 /w:[ 1 3 1 ]
  //: comment g10 @(229,177) /sn:0
  //: /line:"Reset"
  //: /end
  _GGNOR2 #(4) g19 (.I0(w4), .I1(w10), .Z(w8));   //: @(297,219) /sn:0 /w:[ 1 5 5 ]
  //: LED g6 (w8) @(442,204) /sn:0 /w:[ 3 ] /type:0
  //: LED g7 (w10) @(443,346) /sn:0 /w:[ 3 ] /type:0
  _GGNOR2 #(4) g15 (.I0(w8), .I1(w2), .Z(w10));   //: @(315,385) /sn:0 /w:[ 0 0 0 ]
  _GGCLOCK_P100_0_50 g17 (.Z(w6));   //: @(130,426) /sn:0 /w:[ 0 ] /omega:100 /phi:0 /duty:50
  //: joint g5 (w10) @(359, 385) /w:[ 2 4 1 -1 ]
  //: comment g14 @(104,89) /sn:0
  //: /line:"R-S NOR"
  //: /end
  //: SWITCH g0 (w0) @(127,216) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: comment g12 @(444,175) /sn:0
  //: /line:"Q"
  //: /end
  //: joint g18 (w6) @(158, 345) /w:[ 2 4 -1 1 ]

endmodule
//: /netlistEnd

