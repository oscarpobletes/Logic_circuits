//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "bit_adder2.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] B;    //: /sn:0 {0}(#:174,117)(#:174,86){1}
supply0 w7;    //: /sn:0 {0}(539,214)(539,202)(481,202)(481,217){1}
reg [3:0] A;    //: /sn:0 {0}(#:311,82)(311,103){1}
//: {2}(311,104)(311,126){3}
//: {4}(311,127)(311,145){5}
//: {6}(311,146)(311,159){7}
//: {8}(311,160)(311,173){9}
wire w6;    //: /sn:0 {0}(412,378)(412,388)(397,388)(397,347)(390,347)(390,319){1}
wire w16;    //: /sn:0 {0}(231,384)(231,394)(217,394)(217,318){1}
wire w14;    //: /sn:0 {0}(201,218)(201,146)(159,146)(159,123){1}
wire w4;    //: /sn:0 {0}(571,314)(571,344)(501,344)(501,181)(359,181)(359,214)(374,214)(374,219){1}
wire w0;    //: /sn:0 {0}(419,219)(419,127)(315,127){1}
wire w3;    //: /sn:0 {0}(570,384)(570,394)(555,394)(555,314){1}
wire w1;    //: /sn:0 {0}(390,219)(390,140)(179,140)(179,123){1}
wire w8;    //: /sn:0 {0}(322,217)(322,146)(315,146){1}
wire w17;    //: /sn:0 {0}(197,385)(197,395)(212,395)(212,333)(201,333)(201,318){1}
wire a0;    //: /sn:0 {0}(315,104)(323,104)(323,119)(584,119)(584,214){1}
wire b0;    //: /sn:0 {0}(555,214)(555,138)(189,138)(189,123){1}
wire w12;    //: /sn:0 {0}(308,384)(308,394)(293,394)(293,317){1}
wire w11;    //: /sn:0 {0}(309,317)(309,327)(252,327)(252,203)(185,203)(185,218){1}
wire w13;    //: /sn:0 {0}(230,218)(230,160)(306,160){1}
wire w5;    //: /sn:0 {0}(406,319)(406,329)(347,329)(347,202)(277,202)(277,217){1}
wire w9;    //: /sn:0 {0}(293,217)(293,143)(169,143)(169,123){1}
//: enddecls

  //: LED g4 (w12) @(308,377) /sn:0 /w:[ 0 ] /type:0
  adder g8 (.cin(w11), .b(w14), .a(w13), .s(w17), .cout(w16));   //: @(169, 219) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<1 Bo1<1 ]
  assign w13 = A[3]; //: TAP g13 @(309,160) /sn:0 /R:2 /w:[ 1 8 7 ] /ss:0
  //: GROUND g3 (w7) @(481,223) /sn:0 /w:[ 1 ]
  assign w0 = A[1]; //: TAP g2 @(309,127) /sn:0 /R:2 /w:[ 1 4 3 ] /ss:1
  //: LED s0 (w3) @(570,377) /w:[ 0 ] /type:0
  assign a0 = A[0]; //: TAP g1 @(309,104) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  //: comment g16 @(182,18) /sn:0
  //: /line:"4 bits"
  //: /end
  //: DIP g11 (B) @(174,76) /sn:0 /w:[ 1 ] /st:15 /dn:1
  //: DIP g10 (A) @(311,72) /sn:0 /w:[ 0 ] /st:0 /dn:1
  adder g6 (.cin(w4), .b(w1), .a(w0), .s(w6), .cout(w5));   //: @(358, 220) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<1 Bo1<0 ]
  //: LED g9 (w17) @(197,378) /sn:0 /w:[ 0 ] /type:0
  adder g7 (.cin(w5), .b(w9), .a(w8), .s(w12), .cout(w11));   //: @(261, 218) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<1 Bo1<0 ]
  //: LED g15 (w6) @(412,371) /sn:0 /w:[ 0 ] /type:0
  //: LED g5 (w16) @(231,377) /sn:0 /w:[ 0 ] /type:0
  assign {w14, w9, w1, b0} = B; //: CONCAT g14  @(174,118) /sn:0 /R:1 /w:[ 1 1 1 1 0 ] /dr:0 /tp:0 /drp:0
  adder g0 (.a(a0), .b(b0), .cin(w7), .cout(w4), .s(w3));   //: @(523, 215) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>0 Bo0<0 Bo1<1 ]
  assign w8 = A[2]; //: TAP g12 @(309,146) /sn:0 /R:2 /w:[ 1 6 5 ] /ss:1

endmodule
//: /netlistEnd

//: /netlistBegin adder
module adder(cout, s, b, a, cin);
//: interface  /sz:(98, 64) /bd:[ Li0>a(3/64) Li1>b(32/64) Li2>cin(48/64) Ro0<cout(16/64) Ro1<s(32/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input b;    //: /sn:0 {0}(212,44)(78,44)(78,100){1}
//: {2}(76,102)(57,102){3}
//: {4}(78,104)(78,129){5}
//: {6}(80,131)(90,131)(90,132)(131,132){7}
//: {8}(78,133)(78,163)(131,163){9}
input cin;    //: /sn:0 {0}(78,34)(109,34){1}
//: {2}(113,34)(212,34){3}
//: {4}(111,36)(111,96){5}
//: {6}(113,98)(132,98){7}
//: {8}(111,100)(111,127)(131,127){9}
output s;    //: /sn:0 {0}(281,31)(248,31)(248,39)(233,39){1}
input a;    //: /sn:0 {0}(64,69)(87,69){1}
//: {2}(91,69)(199,69)(199,39)(212,39){3}
//: {4}(89,71)(89,81){5}
//: {6}(91,83)(101,83)(101,103)(132,103){7}
//: {8}(89,85)(89,158)(131,158){9}
output cout;    //: /sn:0 {0}(275,106)(228,106){1}
wire w0;    //: /sn:0 {0}(207,101)(153,101){1}
wire w3;    //: /sn:0 {0}(207,111)(167,111)(167,161)(152,161){1}
wire w1;    //: /sn:0 {0}(207,106)(155,106)(155,130)(152,130){1}
//: enddecls

  //: OUT g4 (cout) @(272,106) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g8 (.I0(cin), .I1(b), .Z(w1));   //: @(142,130) /sn:0 /w:[ 9 7 1 ]
  //: OUT g3 (s) @(278,31) /sn:0 /w:[ 0 ]
  //: joint g13 (a) @(89, 83) /w:[ 6 5 -1 8 ]
  //: IN g2 (b) @(55,102) /sn:0 /w:[ 3 ]
  //: IN g1 (a) @(62,69) /sn:0 /w:[ 0 ]
  //: joint g11 (b) @(78, 131) /w:[ 6 5 -1 8 ]
  //: joint g10 (b) @(78, 102) /w:[ -1 1 2 4 ]
  _GGOR3 #(8) g6 (.I0(w0), .I1(w1), .I2(w3), .Z(cout));   //: @(218,106) /sn:0 /w:[ 0 0 0 1 ]
  _GGAND2 #(6) g7 (.I0(cin), .I1(a), .Z(w0));   //: @(143,101) /sn:0 /w:[ 7 7 1 ]
  _GGAND2 #(6) g9 (.I0(a), .I1(b), .Z(w3));   //: @(142,161) /sn:0 /w:[ 9 9 1 ]
  //: joint g15 (cin) @(111, 98) /w:[ 6 5 -1 8 ]
  _GGXOR3 #(11) g5 (.I0(cin), .I1(a), .I2(b), .Z(s));   //: @(223,39) /sn:0 /w:[ 3 3 0 1 ]
  //: joint g14 (cin) @(111, 34) /w:[ 2 -1 1 4 ]
  //: IN g0 (cin) @(76,34) /sn:0 /w:[ 0 ]
  //: joint g12 (a) @(89, 69) /w:[ 2 -1 1 4 ]

endmodule
//: /netlistEnd

