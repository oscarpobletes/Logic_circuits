//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "7_segment_display.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg x1;    //: /sn:0 {0}(487,102)(304,102)(304,132)(294,132){1}
//: {2}(292,130)(292,50)(278,50){3}
//: {4}(292,134)(292,158){5}
//: {6}(294,160)(304,160)(304,161)(420,161){7}
//: {8}(290,160)(280,160)(280,143)(420,143){9}
//: {10}(292,162)(292,179){11}
//: {12}(294,181)(503,181){13}
//: {14}(292,183)(292,212){15}
//: {16}(294,214)(421,214){17}
//: {18}(292,216)(292,235){19}
//: {20}(294,237)(304,237)(304,239)(421,239){21}
//: {22}(292,239)(292,274){23}
//: {24}(294,276)(304,276)(304,273)(421,273){25}
//: {26}(292,278)(292,314){27}
//: {28}(294,316)(304,316)(304,315)(420,315){29}
//: {30}(292,318)(292,348){31}
//: {32}(294,350)(304,350)(304,349)(419,349){33}
//: {34}(292,352)(292,366){35}
//: {36}(294,368)(419,368){37}
//: {38}(292,370)(292,430){39}
//: {40}(294,432)(304,432)(304,421)(421,421){41}
//: {42}(292,434)(292,447){43}
//: {44}(294,449)(304,449)(304,450)(420,450){45}
//: {46}(292,451)(292,470){47}
//: {48}(294,472)(304,472)(304,469)(420,469){49}
//: {50}(292,474)(292,541){51}
reg x0;    //: /sn:0 {0}(503,186)(393,186)(393,188)(383,188){1}
//: {2}(381,186)(381,168){3}
//: {4}(383,166)(420,166){5}
//: {6}(381,164)(381,152){7}
//: {8}(383,150)(393,150)(393,148)(420,148){9}
//: {10}(381,148)(381,95){11}
//: {12}(383,93)(422,93){13}
//: {14}(381,91)(381,53)(357,53){15}
//: {16}(379,93)(369,93)(369,117)(421,117){17}
//: {18}(379,188)(369,188)(369,199)(422,199){19}
//: {20}(381,190)(381,219){21}
//: {22}(383,221)(393,221)(393,219)(421,219){23}
//: {24}(381,223)(381,242){25}
//: {26}(383,244)(421,244){27}
//: {28}(381,246)(381,297){29}
//: {30}(383,299)(393,299)(393,300)(421,300){31}
//: {32}(381,301)(381,320){33}
//: {34}(383,322)(393,322)(393,320)(420,320){35}
//: {36}(381,324)(381,340){37}
//: {38}(383,342)(393,342)(393,344)(419,344){39}
//: {40}(381,344)(381,397){41}
//: {42}(383,399)(393,399)(393,401)(422,401){43}
//: {44}(381,401)(381,444){45}
//: {46}(383,446)(393,446)(393,445)(420,445){47}
//: {48}(381,448)(381,532){49}
reg x3;    //: /sn:0 {0}(507,235)(133,235){1}
//: {2}(131,233)(131,142){3}
//: {4}(133,140)(142,140)(142,107)(487,107){5}
//: {6}(131,138)(131,48)(109,48){7}
//: {8}(131,237)(131,338){9}
//: {10}(133,340)(143,340)(143,361)(514,361){11}
//: {12}(131,342)(131,431){13}
//: {14}(133,433)(143,433)(143,436)(517,436){15}
//: {16}(131,435)(131,535){17}
reg x2;    //: /sn:0 {0}(421,249)(208,249)(208,246)(198,246){1}
//: {2}(196,244)(196,186){3}
//: {4}(198,184)(334,184)(334,156)(483,156){5}
//: {6}(196,182)(196,171){7}
//: {8}(198,169)(208,169)(208,176)(503,176){9}
//: {10}(196,167)(196,116){11}
//: {12}(198,114)(404,114)(404,112)(421,112){13}
//: {14}(196,112)(196,50)(189,50){15}
//: {16}(198,114)(188,114)(188,88)(422,88){17}
//: {18}(198,184)(188,184)(188,194)(422,194){19}
//: {20}(196,248)(196,262){21}
//: {22}(198,264)(208,264)(208,268)(421,268){23}
//: {24}(196,266)(196,297){25}
//: {26}(198,299)(208,299)(208,295)(421,295){27}
//: {28}(196,301)(196,376){29}
//: {30}(198,378)(208,378)(208,373)(419,373){31}
//: {32}(194,378)(184,378)(184,396)(422,396){33}
//: {34}(196,380)(196,416){35}
//: {36}(198,418)(208,418)(208,416)(421,416){37}
//: {38}(196,420)(196,473){39}
//: {40}(198,475)(208,475)(208,474)(420,474){41}
//: {42}(196,477)(196,540){43}
wire w6;    //: /sn:0 {0}(535,368)(615,368)(615,194)(666,194)(666,200){1}
//: {2}(668,202)(681,202)(681,181){3}
//: {4}(666,204)(666,216)(681,216)(681,204){5}
wire w45;    //: /sn:0 {0}(442,419)(489,419)(489,441)(517,441){1}
wire w4;    //: /sn:0 {0}(528,225)(626,225)(626,296)(693,296)(693,279){1}
//: {2}(695,277)(712,277){3}
//: {4}(716,277)(735,277)(735,267){5}
//: {6}(714,275)(714,268){7}
//: {8}(693,275)(693,268){9}
wire w15;    //: /sn:0 {0}(441,146)(483,146){1}
wire w51;    //: /sn:0 {0}(441,472)(502,472)(502,451)(517,451){1}
wire w0;    //: /sn:0 {0}(508,99)(648,99)(648,188)(692,188){1}
//: {2}(696,188)(713,188){3}
//: {4}(717,188)(737,188)(737,162){5}
//: {6}(715,186)(715,176)(716,176)(716,162){7}
//: {8}(694,186)(694,176)(695,176)(695,163){9}
wire w3;    //: /sn:0 {0}(504,151)(591,151)(591,205)(749,205)(749,204){1}
//: {2}(749,200)(749,199){3}
//: {4}(747,202)(735,202)(735,191)(749,191)(749,177){5}
wire w66;    //: /sn:0 {0}(524,181)(584,181)(584,283)(648,283)(648,250)(748,250){1}
//: {2}(750,248)(750,244)(747,244)(747,223){3}
//: {4}(750,252)(750,264)(747,264)(747,244){5}
wire w21;    //: /sn:0 {0}(442,217)(492,217)(492,220)(507,220){1}
wire w76;    //: /sn:0 {0}(516,309)(628,309)(628,270)(671,270){1}
//: {2}(675,270)(681,270)(681,242){3}
//: {4}(673,268)(673,258)(682,258)(682,223){5}
wire w54;    //: /sn:0 {0}(443,399)(499,399)(499,376)(514,376){1}
wire w24;    //: /sn:0 {0}(442,271)(476,271)(476,230)(507,230){1}
wire w36;    //: /sn:0 {0}(440,347)(487,347)(487,366)(514,366){1}
wire w18;    //: /sn:0 {0}(441,164)(459,164)(459,151)(483,151){1}
wire w30;    //: /sn:0 {0}(443,197)(492,197)(492,215)(507,215){1}
wire w12;    //: /sn:0 {0}(442,115)(459,115)(459,97)(487,97){1}
wire w27;    //: /sn:0 {0}(442,244)(466,244)(466,225)(507,225){1}
wire w33;    //: /sn:0 {0}(441,318)(480,318)(480,311)(495,311){1}
wire w48;    //: /sn:0 {0}(441,448)(502,448)(502,446)(517,446){1}
wire w86;    //: /sn:0 {0}(538,443)(602,443)(602,254)(701,254)(701,235){1}
//: {2}(703,233)(722,233)(722,222){3}
//: {4}(701,231)(701,223){5}
wire w9;    //: /sn:0 {0}(443,91)(472,91)(472,92)(487,92){1}
wire w42;    //: /sn:0 {0}(442,298)(480,298)(480,306)(495,306){1}
wire w39;    //: /sn:0 {0}(440,371)(514,371){1}
//: enddecls

  //: LED g4 (w0) @(695,156) /sn:0 /w:[ 9 ] /type:0
  //: joint g8 (w0) @(694, 188) /w:[ 2 8 1 -1 ]
  //: joint g61 (x3) @(131, 140) /w:[ 4 6 -1 3 ]
  //: joint g86 (x2) @(196, 378) /w:[ 30 29 32 34 ]
  //: SWITCH g3 (x3) @(92,48) /sn:0 /w:[ 7 ] /st:0 /dn:1
  //: joint g13 (w66) @(750, 250) /w:[ -1 2 1 4 ]
  //: comment g34 @(630,184) /sn:0
  //: /line:"f"
  //: /end
  _GGAND2 #(6) g37 (.I0(x2), .I1(x0), .Z(w12));   //: @(432,115) /sn:0 /w:[ 13 17 0 ]
  _GGAND2 #(6) g51 (.I0(x2), .I1(!x0), .Z(w54));   //: @(433,399) /sn:0 /w:[ 33 43 0 ]
  _GGOR5 #(12) g55 (.I0(w30), .I1(w21), .I2(w27), .I3(w24), .I4(x3), .Z(w4));   //: @(518,225) /sn:0 /w:[ 1 1 1 1 0 0 ]
  _GGOR4 #(10) g58 (.I0(x3), .I1(w45), .I2(w48), .I3(w51), .Z(w86));   //: @(528,443) /sn:0 /w:[ 15 1 1 1 0 ]
  //: joint g89 (x1) @(292, 449) /w:[ 44 43 -1 46 ]
  //: joint g77 (x3) @(131, 235) /w:[ 1 2 -1 8 ]
  //: joint g76 (x1) @(292, 276) /w:[ 24 23 -1 26 ]
  //: joint g65 (x0) @(381, 166) /w:[ 4 6 -1 3 ]
  //: SWITCH g2 (x2) @(172,50) /sn:0 /w:[ 15 ] /st:0 /dn:1
  //: joint g59 (x0) @(381, 93) /w:[ 12 14 16 11 ]
  //: joint g72 (x1) @(292, 237) /w:[ 20 19 -1 22 ]
  //: SWITCH g1 (x1) @(261,50) /sn:0 /w:[ 3 ] /st:1 /dn:1
  //: joint g64 (x1) @(292, 160) /w:[ 6 5 8 10 ]
  //: LED g11 (w66) @(747,216) /sn:0 /w:[ 3 ] /type:0
  //: LED g16 (w6) @(681,174) /sn:0 /w:[ 3 ] /type:0
  //: joint g87 (x0) @(381, 399) /w:[ 42 41 -1 44 ]
  //: joint g78 (x2) @(196, 299) /w:[ 26 25 -1 28 ]
  //: LED g10 (w3) @(749,192) /sn:0 /w:[ 3 ] /type:0
  //: joint g28 (w6) @(666, 202) /w:[ 2 1 -1 4 ]
  _GGAND2 #(6) g50 (.I0(!x1), .I1(x2), .Z(w51));   //: @(431,472) /sn:0 /w:[ 49 41 0 ]
  //: LED g19 (w66) @(747,237) /sn:0 /w:[ 5 ] /type:0
  //: joint g27 (w86) @(701, 233) /w:[ 2 4 -1 1 ]
  //: comment g32 @(642,301) /sn:0
  //: /line:"d"
  //: /end
  //: joint g69 (x0) @(381, 188) /w:[ 1 2 18 20 ]
  //: LED g6 (w0) @(737,155) /sn:0 /w:[ 5 ] /type:0
  _GGAND2 #(4) g38 (.I0(!x1), .I1(!x0), .Z(w15));   //: @(431,146) /sn:0 /w:[ 9 9 0 ]
  //: joint g75 (x2) @(196, 264) /w:[ 22 21 -1 24 ]
  //: joint g7 (w0) @(715, 188) /w:[ 4 6 3 -1 ]
  //: LED g9 (w3) @(749,170) /sn:0 /w:[ 5 ] /type:0
  _GGOR4 #(10) g57 (.I0(x3), .I1(w36), .I2(w39), .I3(w54), .Z(w6));   //: @(525,368) /sn:0 /w:[ 11 1 1 1 0 ]
  _GGOR3 #(8) g53 (.I0(w15), .I1(w18), .I2(!x2), .Z(w3));   //: @(494,151) /sn:0 /w:[ 1 1 5 0 ]
  //: joint g71 (x0) @(381, 221) /w:[ 22 21 -1 24 ]
  //: LED g20 (w4) @(693,261) /sn:0 /w:[ 9 ] /type:0
  //: LED g15 (w6) @(681,197) /sn:0 /w:[ 5 ] /type:0
  //: comment g31 @(651,276) /sn:0
  //: /line:"c"
  //: /end
  //: joint g68 (x1) @(292, 181) /w:[ 12 11 -1 14 ]
  //: joint g67 (x2) @(196, 169) /w:[ 8 10 -1 7 ]
  _GGAND2 #(6) g39 (.I0(x1), .I1(x0), .Z(w18));   //: @(431,164) /sn:0 /w:[ 7 5 0 ]
  _GGAND2 #(4) g43 (.I0(!x2), .I1(!x0), .Z(w30));   //: @(433,197) /sn:0 /w:[ 19 19 0 ]
  _GGAND2 #(6) g48 (.I0(!x2), .I1(x1), .Z(w45));   //: @(432,419) /sn:0 /w:[ 37 41 0 ]
  //: joint g88 (x0) @(381, 446) /w:[ 46 45 -1 48 ]
  //: joint g73 (x0) @(381, 244) /w:[ 26 25 -1 28 ]
  //: LED g17 (w76) @(682,216) /sn:0 /w:[ 5 ] /type:0
  //: LED g25 (w86) @(701,216) /sn:0 /w:[ 5 ] /type:0
  //: comment g29 @(661,172) /sn:0
  //: /line:"a"
  //: /end
  //: joint g62 (x2) @(196, 114) /w:[ 12 14 16 11 ]
  //: joint g63 (x0) @(381, 150) /w:[ 8 10 -1 7 ]
  _GGAND3 #(8) g42 (.I0(!x1), .I1(x0), .I2(x2), .Z(w27));   //: @(432,244) /sn:0 /w:[ 21 27 0 0 ]
  _GGOR4 #(10) g52 (.I0(w9), .I1(w12), .I2(x1), .I3(x3), .Z(w0));   //: @(498,99) /sn:0 /w:[ 1 1 0 5 0 ]
  //: joint g83 (x0) @(381, 342) /w:[ 38 37 -1 40 ]
  //: joint g74 (x2) @(196, 246) /w:[ 1 2 -1 20 ]
  //: LED g5 (w0) @(716,155) /sn:0 /w:[ 7 ] /type:0
  //: joint g14 (w76) @(673, 270) /w:[ 2 4 1 -1 ]
  _GGOR2 #(6) g56 (.I0(w42), .I1(w33), .Z(w76));   //: @(506,309) /sn:0 /w:[ 1 1 0 ]
  //: joint g94 (x2) @(196, 418) /w:[ 36 35 -1 38 ]
  //: joint g80 (x1) @(292, 316) /w:[ 28 27 -1 30 ]
  //: joint g79 (x0) @(381, 299) /w:[ 30 29 -1 32 ]
  _GGAND2 #(6) g44 (.I0(x1), .I1(!x0), .Z(w33));   //: @(431,318) /sn:0 /w:[ 29 35 0 ]
  _GGAND2 #(4) g47 (.I0(!x2), .I1(!x0), .Z(w42));   //: @(432,298) /sn:0 /w:[ 27 31 0 ]
  //: joint g92 (x3) @(131, 433) /w:[ 14 13 -1 16 ]
  //: joint g85 (x1) @(292, 368) /w:[ 36 35 -1 38 ]
  //: joint g84 (x1) @(292, 350) /w:[ 32 31 -1 34 ]
  //: LED g21 (w4) @(714,261) /sn:0 /w:[ 7 ] /type:0
  //: joint g24 (w4) @(714, 277) /w:[ 4 6 3 -1 ]
  _GGAND2 #(4) g36 (.I0(!x2), .I1(!x0), .Z(w9));   //: @(433,91) /sn:0 /w:[ 17 13 0 ]
  //: joint g23 (w4) @(693, 277) /w:[ 2 8 -1 1 ]
  _GGAND2 #(6) g41 (.I0(!x2), .I1(x1), .Z(w24));   //: @(432,271) /sn:0 /w:[ 23 25 0 ]
  //: joint g93 (x1) @(292, 432) /w:[ 40 39 -1 42 ]
  //: joint g81 (x0) @(381, 322) /w:[ 34 33 -1 36 ]
  _GGAND2 #(6) g40 (.I0(x1), .I1(!x0), .Z(w21));   //: @(432,217) /sn:0 /w:[ 17 23 0 ]
  _GGOR3 #(8) g54 (.I0(x2), .I1(!x1), .I2(x0), .Z(w66));   //: @(514,181) /sn:0 /w:[ 9 13 0 0 ]
  //: joint g60 (x1) @(292, 132) /w:[ 1 2 -1 4 ]
  //: joint g90 (x1) @(292, 472) /w:[ 48 47 -1 50 ]
  //: joint g70 (x1) @(292, 214) /w:[ 16 15 -1 18 ]
  //: SWITCH g0 (x0) @(340,53) /sn:0 /w:[ 15 ] /st:1 /dn:1
  //: LED g22 (w4) @(735,260) /sn:0 /w:[ 5 ] /type:0
  //: LED g26 (w86) @(722,215) /sn:0 /w:[ 3 ] /type:0
  //: comment g35 @(638,241) /sn:0
  //: /line:"g"
  //: /end
  _GGAND2 #(4) g45 (.I0(!x0), .I1(!x1), .Z(w36));   //: @(430,347) /sn:0 /w:[ 39 33 0 ]
  _GGAND2 #(6) g46 (.I0(!x1), .I1(x2), .Z(w39));   //: @(430,371) /sn:0 /w:[ 37 31 0 ]
  //: joint g82 (x3) @(131, 340) /w:[ 10 9 -1 12 ]
  //: joint g66 (x2) @(196, 184) /w:[ 4 6 18 3 ]
  //: LED g18 (w76) @(681,235) /sn:0 /w:[ 3 ] /type:0
  //: joint g12 (w3) @(749, 202) /w:[ -1 2 4 1 ]
  //: joint g91 (x2) @(196, 475) /w:[ 40 39 -1 42 ]
  //: comment g30 @(640,204) /sn:0
  //: /line:"b"
  //: /end
  //: comment g33 @(633,256) /sn:0
  //: /line:"e"
  //: /end
  _GGAND2 #(6) g49 (.I0(!x0), .I1(x1), .Z(w48));   //: @(431,448) /sn:0 /w:[ 47 45 0 ]

endmodule
//: /netlistEnd

