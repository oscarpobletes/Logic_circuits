//: version "2.2"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "Enable.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg x1;    //: /sn:0 {0}(392,95)(417,95)(417,298)(574,298){1}
//: {2}(578,298)(622,298)(622,299)(666,299){3}
//: {4}(576,300)(576,450)(610,450){5}
//: {6}(614,450)(641,450){7}
//: {8}(645,450)(699,450){9}
//: {10}(643,452)(643,601)(729,601){11}
//: {12}(612,452)(612,756)(764,756){13}
supply0 w72;    //: /sn:0 {0}(127,610)(127,573)(331,573){1}
reg x0;    //: /sn:0 {0}(699,434)(685,434){1}
//: {2}(681,434)(671,434){3}
//: {4}(667,434)(634,434)(634,284){5}
//: {6}(636,282)(651,282)(651,283)(666,283){7}
//: {8}(632,282)(627,282)(627,95)(515,95){9}
//: {10}(669,436)(669,585)(729,585){11}
//: {12}(683,436)(683,738)(764,738){13}
supply1 w73;    //: /sn:0 {0}(121,541)(121,557)(331,557){1}
reg x4;    //: /sn:0 {0}(205,677)(291,677)(291,606)(331,606){1}
reg x3;    //: /sn:0 {0}(331,590)(230,590)(230,606)(209,606){1}
reg x2;    //: /sn:0 {0}(270,96)(339,96)(339,314)(491,314){1}
//: {2}(495,314)(580,314)(580,315)(666,315){3}
//: {4}(493,316)(493,466)(544,466){5}
//: {6}(548,466)(597,466){7}
//: {8}(601,466)(699,466){9}
//: {10}(599,468)(599,621)(729,621){11}
//: {12}(546,468)(546,774)(764,774){13}
wire w16;    //: /sn:0 {0}(806,569)(1185,569)(1185,91){1}
wire w6;    //: /sn:0 {0}(841,92)(841,299)(743,299){1}
wire w13;    //: /sn:0 {0}(776,530)(1165,530)(1165,91){1}
wire w65;    //: /sn:0 {0}(442,623)(427,623){1}
wire w7;    //: /sn:0 {0}(873,92)(873,103)(858,103)(858,315)(743,315){1}
wire w50;    //: /sn:0 {0}(806,617)(1247,617)(1247,91){1}
wire w59;    //: /sn:0 {0}(729,673)(522,673)(522,590)(427,590){1}
wire w62;    //: /sn:0 {0}(442,672)(427,672){1}
wire w39;    //: /sn:0 {0}(848,788)(1441,788)(1441,91){1}
wire w4;    //: /sn:0 {0}(778,94)(778,267)(743,267){1}
wire w25;    //: /sn:0 {0}(776,466)(1080,466)(1080,91){1}
wire w56;    //: /sn:0 {0}(848,738)(1378,738)(1378,91){1}
wire w3;    //: /sn:0 {0}(848,809)(1464,809)(1464,91){1}
wire w36;    //: /sn:0 {0}(848,853)(1507,853)(1507,90){1}
wire w22;    //: /sn:0 {0}(806,665)(1316,665)(1316,91){1}
wire w0;    //: /sn:0 {0}(776,418)(1018,418)(1018,91){1}
wire w20;    //: /sn:0 {0}(806,633)(1269,633)(1269,91){1}
wire w30;    //: /sn:0 {0}(776,498)(1122,498)(1122,91){1}
wire w37;    //: /sn:0 {0}(848,828)(1486,828)(1486,90){1}
wire w66;    //: /sn:0 {0}(764,838)(503,838)(503,606)(427,606){1}
wire w18;    //: /sn:0 {0}(806,601)(1227,601)(1227,91){1}
wire w12;    //: /sn:0 {0}(776,482)(1100,482)(1100,91){1}
wire w63;    //: /sn:0 {0}(442,656)(427,656){1}
wire w23;    //: /sn:0 {0}(806,681)(1336,681)(1336,91){1}
wire w10;    //: /sn:0 {0}(961,93)(961,104)(946,104)(946,363)(743,363){1}
wire w21;    //: /sn:0 {0}(806,649)(1290,649)(1290,91){1}
wire w1;    //: /sn:0 {0}(776,434)(1038,434)(1038,91){1}
wire w31;    //: /sn:0 {0}(776,514)(1143,514)(1143,91){1}
wire w68;    //: /sn:0 {0}(427,573)(690,573)(690,523)(699,523){1}
wire w53;    //: /sn:0 {0}(848,720)(1358,720)(1358,91){1}
wire w8;    //: /sn:0 {0}(904,92)(904,103)(889,103)(889,331)(743,331){1}
wire w17;    //: /sn:0 {0}(806,585)(1207,585)(1207,91){1}
wire w69;    //: /sn:0 {0}(427,557)(653,557)(653,373)(666,373){1}
wire w41;    //: /sn:0 {0}(848,756)(1398,756)(1398,91){1}
wire w11;    //: /sn:0 {0}(988,93)(988,379)(743,379){1}
wire w2;    //: /sn:0 {0}(776,450)(1060,450)(1060,91){1}
wire w55;    //: /sn:0 {0}(848,774)(1420,774)(1420,91){1}
wire w5;    //: /sn:0 {0}(807,93)(807,283)(743,283){1}
wire w64;    //: /sn:0 {0}(442,639)(427,639){1}
wire w9;    //: /sn:0 {0}(933,92)(933,103)(918,103)(918,347)(743,347){1}
//: enddecls

  //: joint g44 (x2) @(546, 466) /w:[ 6 -1 5 12 ]
  //: LED g8 (w37) @(1486,83) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g4 (x3) @(192,606) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: SWITCH g3 (x2) @(253,96) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g16 (w0) @(1018,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g26 (w17) @(1207,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g17 (w1) @(1038,84) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g2 (x0) @(498,95) /sn:0 /w:[ 9 ] /st:0 /dn:1
  //: LED g30 (w50) @(1247,84) /sn:0 /w:[ 1 ] /type:0
  DC g23 (.E(w66), .x0(x0), .x1(x1), .x2(x2), .y0(w53), .y1(w56), .y2(w41), .y3(w55), .y4(w39), .y5(w3), .y6(w37), .y7(w36));   //: @(765, 703) /sz:(82, 161) /sn:0 /p:[ Li0>0 Li1>13 Li2>13 Li3>13 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g39 (x2) @(599, 466) /w:[ 8 -1 7 10 ]
  //: LED g24 (w13) @(1165,84) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g1 (x1) @(375,95) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g29 (w18) @(1227,84) /sn:0 /w:[ 1 ] /type:0
  //: LED y4 (w8) @(904,85) /sn:0 /w:[ 0 ] /type:0
  //: LED g18 (w2) @(1060,84) /sn:0 /w:[ 1 ] /type:0
  //: joint g10 (x0) @(669, 434) /w:[ 3 -1 4 10 ]
  //: LED g25 (w16) @(1185,84) /sn:0 /w:[ 1 ] /type:0
  //: LED y0 (w4) @(778,87) /sn:0 /w:[ 0 ] /type:0
  //: LED g6 (w3) @(1464,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g9 (w36) @(1507,83) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g7 (x4) @(188,677) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g35 (w55) @(1420,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g31 (w22) @(1316,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g22 (w31) @(1143,84) /sn:0 /w:[ 1 ] /type:0
  //: GROUND g41 (w72) @(127,616) /sn:0 /w:[ 0 ]
  //: LED g36 (w56) @(1378,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g33 (w53) @(1358,84) /sn:0 /w:[ 1 ] /type:0
  //: joint g40 (x0) @(683, 434) /w:[ 1 -1 2 12 ]
  //: VDD g42 (w73) @(132,541) /sn:0 /w:[ 0 ]
  //: joint g12 (x1) @(643, 450) /w:[ 8 -1 7 10 ]
  //: LED g34 (w39) @(1441,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g28 (w20) @(1269,84) /sn:0 /w:[ 1 ] /type:0
  DC g5 (.x2(x2), .x1(x1), .x0(x0), .E(w59), .y7(w23), .y6(w22), .y5(w21), .y4(w20), .y3(w50), .y2(w18), .y1(w17), .y0(w16));   //: @(730, 553) /sz:(75, 144) /sn:0 /p:[ Li0>11 Li1>11 Li2>11 Li3>0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  DC g11 (.E(w68), .x0(x0), .x1(x1), .x2(x2), .y0(w0), .y1(w1), .y2(w2), .y3(w25), .y4(w12), .y5(w30), .y6(w31), .y7(w13));   //: @(700, 402) /sz:(75, 144) /sn:0 /p:[ Li0>1 Li1>0 Li2>9 Li3>9 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 Ro5<0 Ro6<0 Ro7<0 ]
  //: joint g14 (x1) @(576, 298) /w:[ 2 -1 1 4 ]
  //: LED y1 (w5) @(807,86) /sn:0 /w:[ 0 ] /type:0
  //: LED y2 (w6) @(841,85) /sn:0 /w:[ 0 ] /type:0
  //: LED g19 (w25) @(1080,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g21 (w30) @(1122,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g32 (w23) @(1336,84) /sn:0 /w:[ 1 ] /type:0
  //: LED y3 (w7) @(873,85) /sn:0 /w:[ 0 ] /type:0
  //: LED g20 (w12) @(1100,84) /sn:0 /w:[ 1 ] /type:0
  //: joint g43 (x1) @(612, 450) /w:[ 6 -1 5 12 ]
  DC g38 (.E(w73), .x0(w72), .x1(x3), .x2(x4), .y0(w69), .y1(w68), .y2(w59), .y3(w66), .y4(w65), .y5(w64), .y6(w63), .y7(w62));   //: @(332, 541) /sz:(94, 148) /sn:0 /p:[ Li0>1 Li1>1 Li2>0 Li3>1 Ro0<0 Ro1<0 Ro2<1 Ro3<1 Ro4<1 Ro5<1 Ro6<1 Ro7<1 ]
  DC g0 (.x2(x2), .x1(x1), .x0(x0), .E(w69), .y7(w11), .y6(w10), .y5(w9), .y4(w8), .y3(w7), .y2(w6), .y1(w5), .y0(w4));   //: @(667, 251) /sz:(75, 144) /sn:0 /p:[ Li0>3 Li1>3 Li2>7 Li3>1 Ro0<1 Ro1<1 Ro2<1 Ro3<1 Ro4<1 Ro5<1 Ro6<1 Ro7<1 ]
  //: joint g15 (x2) @(493, 314) /w:[ 2 -1 1 4 ]
  //: LED g27 (w21) @(1290,84) /sn:0 /w:[ 1 ] /type:0
  //: LED g37 (w41) @(1398,84) /sn:0 /w:[ 1 ] /type:0
  //: LED y5 (w9) @(933,85) /sn:0 /w:[ 0 ] /type:0
  //: LED y7 (w11) @(988,86) /sn:0 /w:[ 0 ] /type:0
  //: LED y6 (w10) @(961,86) /sn:0 /w:[ 0 ] /type:0
  //: joint g13 (x0) @(634, 282) /w:[ 6 -1 8 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin DC
module DC(y2, y5, x0, y7, E, y3, y0, x1, y4, y1, y6, x2);
//: interface  /sz:(40, 144) /bd:[ Li0>x2(64/144) Li1>x1(48/144) Li2>x0(32/144) Li3>E(16/144) Ro0<y7(128/144) Ro1<y6(112/144) Ro2<y5(96/144) Ro3<y4(80/144) Ro4<y3(64/144) Ro5<y2(48/144) Ro6<y1(32/144) Ro7<y0(16/144) ] /pd: 0 /pi: 0 /pe: 0 /pp: 1
input x1;    //: /sn:0 {0}(130,-233)(146,-233)(146,-100){1}
//: {2}(148,-98)(160,-98)(160,-96)(272,-96){3}
//: {4}(146,-96)(146,-62){5}
//: {6}(148,-60)(158,-60)(158,-41)(266,-41){7}
//: {8}(146,-58)(146,12){9}
//: {10}(148,14)(158,14)(158,10)(264,10){11}
//: {12}(146,16)(146,66){13}
//: {14}(148,68)(154,68)(154,65)(271,65){15}
//: {16}(146,70)(146,136){17}
//: {18}(148,138)(158,138)(158,128)(271,128){19}
//: {20}(146,140)(146,186){21}
//: {22}(148,188)(158,188)(158,176)(274,176){23}
//: {24}(146,190)(146,223){25}
//: {26}(148,225)(158,225)(158,224)(277,224){27}
//: {28}(146,227)(146,272){29}
//: {30}(148,274)(158,274)(158,269)(277,269){31}
//: {32}(146,276)(146,327){33}
output y4;    //: /sn:0 {0}(383,129)(301,129)(301,130)(292,130){1}
input x0;    //: /sn:0 {0}(66,-224)(74,-224)(74,-99){1}
//: {2}(76,-97)(88,-97)(88,-91)(272,-91){3}
//: {4}(74,-95)(74,-34){5}
//: {6}(76,-32)(86,-32)(86,-36)(266,-36){7}
//: {8}(74,-30)(74,27){9}
//: {10}(76,29)(201,29)(201,15)(264,15){11}
//: {12}(74,31)(74,74){13}
//: {14}(76,76)(86,76)(86,70)(271,70){15}
//: {16}(74,78)(74,152){17}
//: {18}(76,154)(86,154)(86,133)(271,133){19}
//: {20}(74,156)(74,192){21}
//: {22}(76,194)(86,194)(86,181)(274,181){23}
//: {24}(74,196)(74,230){25}
//: {26}(76,232)(84,232)(84,229)(277,229){27}
//: {28}(74,234)(74,286){29}
//: {30}(76,288)(85,288)(85,317)(125,317)(125,295)(175,295)(175,274)(277,274){31}
//: {32}(74,290)(74,339){33}
output y0;    //: /sn:0 {0}(378,-96)(308,-96)(308,-94)(293,-94){1}
output y1;    //: /sn:0 {0}(383,-41)(302,-41)(302,-39)(287,-39){1}
output y2;    //: /sn:0 {0}(385,3)(300,3)(300,12)(285,12){1}
output y3;    //: /sn:0 {0}(380,64)(307,64)(307,67)(292,67){1}
input E;    //: /sn:0 {0}(-20,349)(241,349)(241,283){1}
//: {2}(243,281)(253,281)(253,279)(277,279){3}
//: {4}(241,279)(241,233){5}
//: {6}(243,231)(253,231)(253,234)(277,234){7}
//: {8}(241,229)(241,187){9}
//: {10}(243,185)(253,185)(253,186)(274,186){11}
//: {12}(241,183)(241,140){13}
//: {14}(243,138)(271,138){15}
//: {16}(241,136)(241,77){17}
//: {18}(243,75)(271,75){19}
//: {20}(241,73)(241,22){21}
//: {22}(243,20)(264,20){23}
//: {24}(241,18)(241,-29){25}
//: {26}(243,-31)(266,-31){27}
//: {28}(241,-33)(241,-86)(272,-86){29}
output y5;    //: /sn:0 {0}(401,174)(310,174)(310,178)(295,178){1}
output y7;    //: /sn:0 {0}(391,274)(313,274)(313,271)(298,271){1}
input x2;    //: /sn:0 {0}(210,-225)(221,-225)(221,-104){1}
//: {2}(223,-102)(235,-102)(235,-101)(272,-101){3}
//: {4}(221,-100)(221,-47){5}
//: {6}(223,-45)(233,-45)(233,-46)(266,-46){7}
//: {8}(221,-43)(221,-17){9}
//: {10}(223,-15)(229,-15)(229,5)(264,5){11}
//: {12}(221,-13)(221,53){13}
//: {14}(223,55)(233,55)(233,60)(271,60){15}
//: {16}(221,57)(221,118){17}
//: {18}(223,120)(233,120)(233,123)(271,123){19}
//: {20}(221,122)(221,170){21}
//: {22}(223,172)(233,172)(233,171)(274,171){23}
//: {24}(221,174)(221,219){25}
//: {26}(223,221)(233,221)(233,219)(277,219){27}
//: {28}(221,223)(221,258){29}
//: {30}(223,260)(233,260)(233,264)(277,264){31}
//: {32}(221,262)(221,333){33}
output y6;    //: /sn:0 {0}(393,228)(314,228)(314,226)(298,226){1}
//: enddecls

  _GGAND4 #(10) g4 (.I0(!x2), .I1(!x1), .I2(x0), .I3(E), .Z(y4));   //: @(282,130) /sn:0 /w:[ 19 19 19 15 1 ]
  //: OUT g44 (y2) @(382,3) /sn:0 /w:[ 0 ]
  //: joint g8 (x2) @(221, -102) /w:[ 2 1 -1 4 ]
  _GGAND4 #(10) g3 (.I0(x2), .I1(x1), .I2(!x0), .I3(E), .Z(y3));   //: @(282,67) /sn:0 /w:[ 15 15 15 19 1 ]
  //: joint g16 (x1) @(146, -60) /w:[ 6 5 -1 8 ]
  //: OUT g47 (y5) @(398,174) /sn:0 /w:[ 0 ]
  //: joint g17 (x1) @(146, 14) /w:[ 10 9 -1 12 ]
  //: joint g26 (x2) @(221, 172) /w:[ 22 21 -1 24 ]
  _GGAND4 #(10) g2 (.I0(!x2), .I1(x1), .I2(!x0), .I3(E), .Z(y2));   //: @(275,12) /sn:0 /w:[ 11 11 11 23 1 ]
  //: joint g23 (x1) @(146, 138) /w:[ 18 17 -1 20 ]
  //: joint g30 (x1) @(146, 225) /w:[ 26 25 -1 28 ]
  _GGAND4 #(10) g1 (.I0(x2), .I1(!x1), .I2(!x0), .I3(E), .Z(y1));   //: @(277,-39) /sn:0 /w:[ 7 7 7 27 1 ]
  //: joint g24 (x2) @(221, 120) /w:[ 18 17 -1 20 ]
  //: joint g39 (E) @(241, 185) /w:[ 10 12 -1 9 ]
  //: joint g29 (x0) @(74, 232) /w:[ 26 25 -1 28 ]
  //: IN g51 (x0) @(64,-224) /sn:0 /w:[ 0 ]
  //: joint g18 (x2) @(221, -15) /w:[ 10 9 -1 12 ]
  //: joint g25 (x0) @(74, 154) /w:[ 18 17 -1 20 ]
  //: OUT g49 (y7) @(388,274) /sn:0 /w:[ 0 ]
  _GGAND4 #(10) g6 (.I0(x2), .I1(!x1), .I2(x0), .I3(E), .Z(y5));   //: @(285,178) /sn:0 /w:[ 23 23 23 11 1 ]
  //: IN g50 (E) @(-22,349) /sn:0 /w:[ 0 ]
  _GGAND4 #(10) g7 (.I0(!x2), .I1(x1), .I2(x0), .I3(E), .Z(y6));   //: @(288,226) /sn:0 /w:[ 27 27 27 7 1 ]
  //: joint g35 (E) @(241, 20) /w:[ 22 24 -1 21 ]
  //: joint g22 (x0) @(74, 76) /w:[ 14 13 -1 16 ]
  //: joint g31 (x2) @(221, 260) /w:[ 30 29 -1 32 ]
  //: joint g36 (E) @(241, 75) /w:[ 18 20 -1 17 ]
  //: joint g41 (E) @(241, 281) /w:[ 2 4 -1 1 ]
  //: OUT g45 (y3) @(377,64) /sn:0 /w:[ 0 ]
  //: joint g33 (x0) @(74, 288) /w:[ 30 29 -1 32 ]
  //: joint g40 (E) @(241, 231) /w:[ 6 8 -1 5 ]
  //: OUT g42 (y0) @(375,-96) /sn:0 /w:[ 0 ]
  //: IN g52 (x1) @(128,-233) /sn:0 /w:[ 0 ]
  //: joint g12 (x0) @(74, -97) /w:[ 2 1 -1 4 ]
  //: joint g28 (x2) @(221, 221) /w:[ 26 25 -1 28 ]
  //: joint g34 (E) @(241, -31) /w:[ 26 28 -1 25 ]
  //: OUT g46 (y4) @(380,129) /sn:0 /w:[ 0 ]
  _GGAND4 #(10) g5 (.I0(x2), .I1(x1), .I2(x0), .I3(E), .Z(y7));   //: @(288,271) /sn:0 /w:[ 31 31 31 3 1 ]
  //: joint g14 (x2) @(221, -45) /w:[ 6 5 -1 8 ]
  //: joint g19 (x0) @(74, 29) /w:[ 10 9 -1 12 ]
  //: joint g21 (x1) @(146, 68) /w:[ 14 13 -1 16 ]
  //: joint g20 (x2) @(221, 55) /w:[ 14 13 -1 16 ]
  //: joint g32 (x1) @(146, 274) /w:[ 30 29 -1 32 ]
  _GGAND4 #(10) g0 (.I0(!x2), .I1(!x1), .I2(!x0), .I3(E), .Z(y0));   //: @(283,-94) /sn:0 /w:[ 3 3 3 29 1 ]
  //: joint g15 (x0) @(74, -32) /w:[ 6 5 -1 8 ]
  //: joint g38 (x0) @(74, 194) /w:[ 22 21 -1 24 ]
  //: OUT g43 (y1) @(380,-41) /sn:0 /w:[ 0 ]
  //: joint g27 (x1) @(146, 188) /w:[ 22 21 -1 24 ]
  //: OUT g48 (y6) @(390,228) /sn:0 /w:[ 0 ]
  //: joint g37 (E) @(241, 138) /w:[ 14 16 -1 13 ]
  //: IN g53 (x2) @(208,-225) /sn:0 /w:[ 0 ]
  //: joint g13 (x1) @(146, -98) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

