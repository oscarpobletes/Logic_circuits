//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg x1;    //: /sn:0 {0}(239,263)(266,263)(266,299){1}
//: {2}(268,301)(428,301){3}
//: {4}(266,303)(266,350){5}
//: {6}(268,352)(351,352)(351,355)(422,355){7}
//: {8}(266,354)(266,402){9}
//: {10}(268,404)(278,404)(278,402)(424,402){11}
//: {12}(266,406)(266,453){13}
//: {14}(268,455)(278,455)(278,454)(427,454){15}
//: {16}(266,457)(266,510){17}
//: {18}(268,512)(278,512)(278,506)(431,506){19}
//: {20}(266,514)(266,578){21}
reg x0;    //: /sn:0 {0}(431,511)(361,511)(361,517)(351,517){1}
//: {2}(349,515)(349,460){3}
//: {4}(351,458)(361,458)(361,459)(427,459){5}
//: {6}(349,456)(349,409){7}
//: {8}(351,407)(424,407){9}
//: {10}(349,405)(349,365){11}
//: {12}(351,363)(361,363)(361,360)(422,360){13}
//: {14}(349,361)(349,314){15}
//: {16}(351,312)(361,312)(361,311)(428,311){17}
//: {18}(349,310)(349,263)(325,263){19}
//: {20}(349,519)(349,568){21}
reg x2;    //: /sn:0 {0}(428,291)(163,291){1}
//: {2}(161,289)(161,260)(146,260){3}
//: {4}(161,293)(161,349){5}
//: {6}(163,351)(173,351)(173,350)(422,350){7}
//: {8}(161,353)(161,387){9}
//: {10}(163,389)(173,389)(173,397)(424,397){11}
//: {12}(161,391)(161,444){13}
//: {14}(163,446)(173,446)(173,449)(427,449){15}
//: {16}(161,448)(161,501){17}
//: {18}(163,503)(173,503)(173,501)(431,501){19}
//: {20}(161,505)(161,575){21}
wire w16;    //: /sn:0 {0}(467,401)(467,417)(535,417){1}
wire w14;    //: /sn:0 {0}(535,427)(476,427)(476,506)(452,506){1}
wire [2:0] w21;    //: /sn:0 {0}(#:434,301)(498,301){1}
//: {2}(#:502,301)(600,301)(600,285){3}
//: {4}(500,299)(500,283){5}
wire w18;    //: /sn:0 {0}(535,422)(471,422)(471,454){1}
wire w8;    //: /sn:0 {0}(445,402)(460,402){1}
wire w11;    //: /sn:0 {0}(448,454)(463,454){1}
wire w5;    //: /sn:0 {0}(443,355)(520,355)(520,412)(535,412){1}
wire Y;    //: /sn:0 {0}(631,404)(631,419)(556,419){1}
//: enddecls

  _GGOR4 #(10) g8 (.I0(w5), .I1(w16), .I2(w18), .I3(w14), .Z(Y));   //: @(546,419) /sn:0 /w:[ 1 1 0 0 1 ]
  _GGAND3 #(8) g4 (.I0(!x2), .I1(x1), .I2(x0), .Z(w5));   //: @(433,355) /sn:0 /w:[ 7 7 13 0 ]
  //: joint g13 (x2) @(161, 291) /w:[ 1 2 -1 4 ]
  //: comment g3 @(115,68) /sn:0
  //: /line:"Given three bits indicate when the majority are 1"
  //: /line:""
  //: /line:"x2 x1 x0 | Majority ones"
  //: /line:"0  0   0       0"
  //: /line:"0  0   1       0"
  //: /line:"0  1   0       0"
  //: /line:"0  1   1       1"
  //: /line:"1  0   0       0"
  //: /line:"1  0   1       1"
  //: /line:"1  1   0       1"
  //: /line:"1  1   1       1"
  //: /end
  //: SWITCH g2 (x0) @(308,263) /sn:0 /w:[ 19 ] /st:0 /dn:1
  //: SWITCH g1 (x1) @(222,263) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g16 (w21) @(500, 301) /w:[ 2 4 1 -1 ]
  //: LED g11 (w21) @(600,278) /sn:0 /w:[ 3 ] /type:3
  //: comment g28 @(504,322) /sn:0
  //: /line:"3 bits bus"
  //: /line:""
  //: /end
  //: LED g10 (w21) @(500,276) /sn:0 /w:[ 5 ] /type:1
  //: joint g27 (x0) @(349, 517) /w:[ 1 2 -1 20 ]
  //: joint g19 (x2) @(161, 389) /w:[ 10 9 -1 12 ]
  _GGAND3 #(8) g6 (.I0(x2), .I1(x1), .I2(!x0), .Z(w11));   //: @(438,454) /sn:0 /w:[ 15 15 5 0 ]
  //: joint g9 (x2) @(161, 351) /w:[ 6 5 -1 8 ]
  _GGAND3 #(8) g7 (.I0(x2), .I1(x1), .I2(x0), .Z(w14));   //: @(442,506) /sn:0 /w:[ 19 19 0 1 ]
  //: joint g20 (x1) @(266, 404) /w:[ 10 9 -1 12 ]
  //: joint g15 (x0) @(349, 312) /w:[ 16 18 -1 15 ]
  //: comment g29 @(661,403) /sn:0
  //: /line:"Most ones?"
  //: /end
  //: joint g25 (x2) @(161, 503) /w:[ 18 17 -1 20 ]
  //: joint g17 (x1) @(266, 352) /w:[ 6 5 -1 8 ]
  //: joint g14 (x1) @(266, 301) /w:[ 2 1 -1 4 ]
  _GGAND3 #(8) g5 (.I0(x2), .I1(!x1), .I2(x0), .Z(w8));   //: @(435,402) /sn:0 /w:[ 11 11 9 0 ]
  //: joint g24 (x0) @(349, 458) /w:[ 4 6 -1 3 ]
  //: joint g21 (x0) @(349, 407) /w:[ 8 10 -1 7 ]
  //: joint g23 (x1) @(266, 455) /w:[ 14 13 -1 16 ]
  //: joint g26 (x1) @(266, 512) /w:[ 18 17 -1 20 ]
  //: joint g22 (x2) @(161, 446) /w:[ 14 13 -1 16 ]
  //: SWITCH g0 (x2) @(129,260) /sn:0 /w:[ 3 ] /st:0 /dn:1
  //: joint g18 (x0) @(349, 363) /w:[ 12 14 -1 11 ]
  assign w21 = {x2, x1, x0}; //: CONCAT g12  @(433,301) /sn:0 /w:[ 0 0 3 17 ] /dr:0 /tp:0 /drp:1
  //: LED Y (Y) @(631,397) /w:[ 0 ] /type:0

endmodule
//: /netlistEnd

