//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
output Q;    //: /sn:0 {0}(541,100)(485,100)(485,106)(470,106){1}
output notQ;    //: /sn:0 {0}(470,122)(510,122)(510,128)(531,128){1}
input Clk;    //: /sn:0 {0}(79,144)(138,144)(138,156)(153,156){1}
input notE;    //: /sn:0 {0}(81,185)(140,185)(140,161)(153,161){1}
input D;    //: /sn:0 {0}(237,146)(171,146)(171,128)(102,128)(102,106){1}
//: {2}(104,104)(114,104)(114,95)(237,95){3}
//: {4}(102,102)(102,92)(70,92){5}
wire w1;    //: /sn:0 {0}(174,159)(196,159){1}
//: {2}(200,159)(224,159)(224,151)(237,151){3}
//: {4}(198,157)(198,100)(237,100){5}
wire w2;    //: /sn:0 {0}(258,98)(285,98)(285,122)(335,122){1}
wire w5;    //: /sn:0 {0}(258,149)(302,149)(302,106)(335,106){1}
//: enddecls

  RS_trigger g8 (.R(w5), .S(w2), .notQ(Q), .Q(notQ));   //: @(336, 90) /sz:(133, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<0 ]
  _GGAND2 #(6) g4 (.I0(!D), .I1(w1), .Z(w5));   //: @(248,149) /sn:0 /w:[ 0 3 0 ]
  _GGAND2 #(6) g3 (.I0(D), .I1(w1), .Z(w2));   //: @(248,98) /sn:0 /w:[ 3 5 0 ]
  //: IN g2 (notE) @(79,185) /sn:0 /w:[ 0 ]
  //: IN g1 (Clk) @(77,144) /sn:0 /w:[ 0 ]
  //: OUT g10 (notQ) @(528,128) /sn:0 /w:[ 1 ]
  //: joint g6 (D) @(102, 104) /w:[ 2 4 -1 1 ]
  //: OUT g9 (Q) @(538,100) /sn:0 /w:[ 0 ]
  //: joint g7 (w1) @(198, 159) /w:[ 2 4 1 -1 ]
  _GGAND2 #(6) g5 (.I0(Clk), .I1(!notE), .Z(w1));   //: @(164,159) /sn:0 /w:[ 1 1 0 ]
  //: IN g0 (D) @(68,92) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin RS_trigger
module RS_trigger(Q, R, notQ, S);
//: interface  /sz:(133, 48) /bd:[ Li0>S(32/48) Li1>R(16/48) Ro0<Q(32/48) Ro1<notQ(16/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Q;    //: /sn:0 {0}(471,118)(450,118)(450,119)(326,119){1}
//: {2}(322,119)(264,119){3}
//: {4}(324,121)(324,187)(230,187)(230,202)(240,202){5}
output notQ;    //: /sn:0 {0}(465,200)(306,200){1}
//: {2}(304,198)(304,136)(233,136)(233,121)(243,121){3}
//: {4}(302,200)(261,200){5}
input R;    //: /sn:0 {0}(240,197)(102,197)(102,207)(74,207){1}
input S;    //: /sn:0 {0}(73,134)(188,134)(188,116)(243,116){1}
//: enddecls

  //: OUT g4 (Q) @(468,118) /sn:0 /w:[ 0 ]
  _GGNAND2 #(4) g3 (.I0(R), .I1(Q), .Z(notQ));   //: @(251,200) /sn:0 /w:[ 0 5 5 ]
  _GGNAND2 #(4) g2 (.I0(S), .I1(notQ), .Z(Q));   //: @(254,119) /sn:0 /w:[ 1 3 3 ]
  //: IN g1 (R) @(72,207) /sn:0 /w:[ 1 ]
  //: joint g6 (Q) @(324, 119) /w:[ 1 -1 2 4 ]
  //: joint g7 (notQ) @(304, 200) /w:[ 1 2 4 -1 ]
  //: OUT g5 (notQ) @(462,200) /sn:0 /w:[ 0 ]
  //: IN g0 (S) @(71,134) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

