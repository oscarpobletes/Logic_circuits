//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "substraction_using_addition_8bits.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] w6;    //: /sn:0 {0}(#:246,116)(246,147){1}
//: {2}(#:248,149)(663,149)(663,93){3}
//: {4}(246,151)(246,231)(345,231)(345,244){5}
reg [7:0] w7;    //: /sn:0 {0}(#:391,123)(391,147)(390,147)(390,151){1}
//: {2}(#:392,153)(517,153)(517,94){3}
//: {4}(390,155)(390,234)(377,234)(377,244){5}
supply0 w5;    //: /sn:0 {0}(283,351)(283,325)(200,325)(200,330){1}
supply1 w9;    //: /sn:0 {0}(385,258)(405,258)(405,316)(430,316)(430,338){1}
//: {2}(432,340)(473,340)(473,303){3}
//: {4}(430,342)(430,365)(323,365){5}
wire w14;    //: /sn:0 {0}(557,259)(557,388)(336,388)(336,476)(350,476){1}
//: {2}(354,476)(368,476){3}
//: {4}(352,474)(352,338){5}
//: {6}(352,478)(352,528)(412,528)(412,538)(429,538){7}
wire w4;    //: /sn:0 {0}(337,258)(322,258){1}
wire [7:0] w15;    //: /sn:0 {0}(468,462)(448,462)(#:448,451)(#:433,451){1}
wire w3;    //: /sn:0 {0}(257,365)(275,365){1}
wire [7:0] w21;    //: /sn:0 {0}(#:299,380)(299,533)(#:429,533){1}
wire [7:0] w1;    //: /sn:0 {0}(#:489,465)(613,465)(#:613,268){1}
wire w8;    //: /sn:0 {0}(384,476)(405,476)(405,453)(412,453){1}
wire [7:0] w18;    //: /sn:0 {0}(468,467)(465,467)(#:465,536)(#:450,536){1}
wire [7:0] w2;    //: /sn:0 {0}(#:412,448)(382,448)(382,322)(365,322)(365,334)(352,334){1}
//: {2}(351,334)(339,334)(339,293){3}
//: {4}(341,291)(361,291)(#:361,273){5}
//: {6}(337,291)(315,291)(315,351){7}
//: enddecls

  _GGNBUF #(2) g4 (.I(w14), .Z(w8));   //: @(374,476) /sn:0 /w:[ 3 0 ]
  //: LED g8 (w14) @(557,252) /sn:0 /w:[ 0 ] /type:0
  //: DIP g3 (w7) @(391,113) /sn:0 /w:[ 0 ] /st:6 /dn:1
  //: DIP g2 (w6) @(246,106) /sn:0 /w:[ 0 ] /st:4 /dn:1
  //: LED g1 (w1) @(613,261) /sn:0 /w:[ 1 ] /type:3
  //: VDD g11 (w9) @(484,303) /sn:0 /w:[ 3 ]
  //: GROUND g16 (w5) @(200,336) /sn:0 /w:[ 1 ]
  _GGAND2x8 #(6) g10 (.I0(w2), .I1({8{w8}}), .Z(w15));   //: @(423,451) /sn:0 /w:[ 0 1 1 ]
  //: joint g6 (w2) @(339, 291) /w:[ 4 -1 6 3 ]
  //: joint g7 (w14) @(352, 476) /w:[ 2 4 1 6 ]
  _GGOR2x8 #(6) g9 (.I0(w15), .I1(w18), .Z(w1));   //: @(479,465) /sn:0 /w:[ 0 0 0 ]
  //: comment g15 @(515,197) /sn:0
  //: /line:"Most significant bit (-)"
  //: /line:"          |"
  //: /line:"          v"
  //: /end
  assign w14 = w2[0]; //: TAP g17 @(352,332) /sn:0 /R:1 /w:[ 5 2 1 ] /ss:1
  //: joint g25 (w7) @(390, 153) /w:[ 2 1 -1 4 ]
  _GGADD8 #(70, 72, 62, 64) g5 (.A(w5), .B(~w2), .S(w21), .CI(w9), .CO(w3));   //: @(299,367) /sn:0 /w:[ 0 7 0 5 1 ]
  _GGAND2x8 #(6) g14 (.I0(w21), .I1({8{w14}}), .Z(w18));   //: @(440,536) /sn:0 /w:[ 1 7 1 ]
  //: comment g21 @(564,159) /sn:0
  //: /line:"-------"
  //: /line:"-------"
  //: /end
  //: joint g24 (w6) @(246, 149) /w:[ 2 1 -1 4 ]
  //: LED g23 (w7) @(517,87) /sn:0 /w:[ 3 ] /type:3
  _GGADD8 #(70, 72, 62, 64) g0 (.A(~w6), .B(w7), .S(w2), .CI(w9), .CO(w4));   //: @(361,260) /sn:0 /w:[ 5 5 5 0 0 ]
  //: LED g22 (w6) @(663,86) /sn:0 /w:[ 3 ] /type:3
  //: comment g26 @(572,70) /sn:0
  //: /line:"------"
  //: /line:""
  //: /end
  //: joint g12 (w9) @(430, 340) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

