//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "nums.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [3:0] w0;    //: /sn:0 {0}(#:210,115)(#:210,87){1}
wire w32;    //: /sn:0 {0}(985,81)(985,102)(854,102)(854,334)(594,334){1}
wire w6;    //: /sn:0 {0}(521,354)(491,354)(491,596)(463,596){1}
wire w7;    //: /sn:0 {0}(374,153)(425,153)(425,196)(440,196){1}
wire w14;    //: /sn:0 {0}(521,304)(483,304)(483,206)(461,206){1}
wire w16;    //: /sn:0 {0}(440,206)(376,206){1}
wire w19;    //: /sn:0 {0}(884,127)(884,140){1}
//: {2}(886,142)(899,142){3}
//: {4}(903,142)(915,142){5}
//: {6}(919,142)(931,142){7}
//: {8}(935,142)(947,142){9}
//: {10}(951,142)(963,142){11}
//: {12}(967,142)(979,142){13}
//: {14}(983,142)(997,142)(997,127){15}
//: {16}(981,140)(981,127){17}
//: {18}(965,140)(965,127){19}
//: {20}(949,140)(949,127){21}
//: {22}(933,140)(933,127){23}
//: {24}(917,140)(917,127){25}
//: {26}(901,140)(901,127){27}
//: {28}(884,144)(884,344)(594,344){29}
wire w4;    //: /sn:0 {0}(594,324)(850,324)(850,101)(902,101)(902,81){1}
wire w15;    //: /sn:0 {0}(521,364)(500,364)(500,641)(438,641){1}
wire w3;    //: /sn:0 {0}(887,197)(887,203)(654,203)(654,413){1}
//: {2}(656,415)(669,415){3}
//: {4}(673,415)(685,415){5}
//: {6}(689,415)(701,415){7}
//: {8}(705,415)(717,415){9}
//: {10}(721,415)(733,415){11}
//: {12}(737,415)(749,415){13}
//: {14}(753,415)(1000,415)(1000,197){15}
//: {16}(751,413)(751,203)(984,203)(984,197){17}
//: {18}(735,413)(735,203)(968,203)(968,197){19}
//: {20}(719,413)(719,203)(952,203)(952,197){21}
//: {22}(703,413)(703,203)(936,203)(936,197){23}
//: {24}(687,413)(687,203)(920,203)(920,197){25}
//: {26}(671,413)(671,203)(904,203)(904,197){27}
//: {28}(652,415)(635,415)(635,364)(594,364){29}
wire w34;    //: /sn:0 {0}(417,649)(327,649){1}
//: {2}(325,647)(325,539){3}
//: {4}(327,537)(354,537){5}
//: {6}(325,535)(325,493){7}
//: {8}(327,491)(377,491){9}
//: {10}(325,489)(325,463){11}
//: {12}(327,461)(350,461){13}
//: {14}(325,459)(325,430){15}
//: {16}(327,428)(376,428){17}
//: {18}(325,426)(325,403){19}
//: {20}(327,401)(348,401){21}
//: {22}(325,399)(325,389){23}
//: {24}(327,387)(376,387){25}
//: {26}(325,385)(325,361){27}
//: {28}(327,359)(347,359){29}
//: {30}(325,357)(325,335){31}
//: {32}(327,333)(376,333){33}
//: {34}(325,331)(325,304){35}
//: {36}(327,302)(347,302){37}
//: {38}(325,300)(325,267){39}
//: {40}(327,265)(355,265){41}
//: {42}(325,263)(325,243){43}
//: {44}(327,241)(377,241){45}
//: {46}(325,239)(325,213){47}
//: {48}(327,211)(355,211){49}
//: {50}(325,209)(325,186){51}
//: {52}(327,184)(375,184){53}
//: {54}(325,182)(325,152){55}
//: {56}(327,150)(353,150){57}
//: {58}(325,148)(325,134)(225,134)(225,121){59}
//: {60}(325,651)(325,681)(391,681){61}
wire w75;    //: /sn:0 {0}(521,324)(491,324)(491,316){1}
//: {2}(493,314)(521,314){3}
//: {4}(489,314)(460,314){5}
wire w76;    //: /sn:0 {0}(521,334)(475,334)(475,462)(459,462){1}
wire w21;    //: /sn:0 {0}(397,328)(413,328)(413,312)(439,312){1}
wire w31;    //: /sn:0 {0}(394,604)(427,604)(427,598)(442,598){1}
wire w28;    //: /sn:0 {0}(885,164)(885,170)(653,170)(653,368){1}
//: {2}(655,370)(668,370){3}
//: {4}(672,370)(684,370){5}
//: {6}(688,370)(700,370){7}
//: {8}(704,370)(716,370){9}
//: {10}(720,370)(732,370){11}
//: {12}(736,370)(748,370){13}
//: {14}(752,370)(998,370)(998,164){15}
//: {16}(750,368)(750,170)(982,170)(982,164){17}
//: {18}(734,368)(734,170)(966,170)(966,164){19}
//: {20}(718,368)(718,170)(950,170)(950,164){21}
//: {22}(702,368)(702,170)(934,170)(934,164){23}
//: {24}(686,368)(686,170)(918,170)(918,164){25}
//: {26}(670,368)(670,170)(902,170)(902,164){27}
//: {28}(651,370)(642,370)(642,354)(594,354){29}
wire w20;    //: /sn:0 {0}(440,211)(413,211)(413,233)(398,233){1}
wire w23;    //: /sn:0 {0}(440,216)(420,216)(420,257)(376,257){1}
wire w24;    //: /sn:0 {0}(442,593)(387,593)(387,578)(372,578){1}
wire w36;    //: /sn:0 {0}(521,374)(509,374)(509,673)(412,673){1}
wire [7:0] w1;    //: /sn:0 {0}(#:588,339)(#:527,339){1}
wire w25;    //: /sn:0 {0}(439,317)(419,317)(419,351)(368,351){1}
wire w18;    //: /sn:0 {0}(438,462)(404,462)(404,468)(371,468){1}
wire w35;    //: /sn:0 {0}(594,304)(841,304)(841,99)(932,99)(932,81){1}
wire w8;    //: /sn:0 {0}(396,283)(424,283)(424,302)(439,302){1}
wire w30;    //: /sn:0 {0}(417,644)(243,644){1}
//: {2}(241,642)(241,608){3}
//: {4}(243,606)(373,606){5}
//: {6}(241,604)(241,561){7}
//: {8}(243,559)(381,559){9}
//: {10}(241,557)(241,498){11}
//: {12}(243,496)(377,496){13}
//: {14}(241,494)(241,468){15}
//: {16}(243,466)(350,466){17}
//: {18}(241,464)(241,435){19}
//: {20}(243,433)(376,433){21}
//: {22}(241,431)(241,408){23}
//: {24}(243,406)(348,406){25}
//: {26}(241,404)(241,384){27}
//: {28}(243,382)(376,382){29}
//: {30}(241,380)(241,356){31}
//: {32}(243,354)(347,354){33}
//: {34}(241,352)(241,330){35}
//: {36}(243,328)(376,328){37}
//: {38}(241,326)(241,314){39}
//: {40}(243,312)(347,312){41}
//: {42}(241,310)(241,290){43}
//: {44}(243,288)(375,288){45}
//: {46}(241,286)(241,262){47}
//: {48}(243,260)(355,260){49}
//: {50}(241,258)(241,238){51}
//: {52}(243,236)(377,236){53}
//: {54}(241,234)(241,181){55}
//: {56}(243,179)(375,179){57}
//: {58}(241,177)(241,145)(215,145)(215,121){59}
//: {60}(241,646)(241,676)(391,676){61}
wire w17;    //: /sn:0 {0}(439,531)(417,531)(417,557)(402,557){1}
wire w22;    //: /sn:0 {0}(353,155)(166,155){1}
//: {2}(164,153)(164,143)(205,143)(205,121){3}
//: {4}(164,157)(164,172){5}
//: {6}(166,174)(375,174){7}
//: {8}(164,176)(164,204){9}
//: {10}(166,206)(355,206){11}
//: {12}(164,208)(164,229){13}
//: {14}(166,231)(377,231){15}
//: {16}(164,233)(164,253){17}
//: {18}(166,255)(355,255){19}
//: {20}(164,257)(164,281){21}
//: {22}(166,283)(375,283){23}
//: {24}(164,285)(164,321){25}
//: {26}(166,323)(376,323){27}
//: {28}(164,325)(164,347){29}
//: {30}(166,349)(347,349){31}
//: {32}(164,351)(164,375){33}
//: {34}(166,377)(376,377){35}
//: {36}(164,379)(164,409){37}
//: {38}(166,411)(348,411){39}
//: {40}(164,413)(164,436){41}
//: {42}(166,438)(376,438){43}
//: {44}(164,440)(164,469){45}
//: {46}(166,471)(350,471){47}
//: {48}(164,473)(164,499){49}
//: {50}(166,501)(377,501){51}
//: {52}(164,503)(164,530){53}
//: {54}(166,532)(354,532){55}
//: {56}(164,534)(164,552){57}
//: {58}(166,554)(381,554){59}
//: {60}(164,556)(164,578){61}
//: {62}(166,580)(351,580){63}
//: {64}(164,582)(164,637){65}
//: {66}(166,639)(417,639){67}
//: {68}(164,641)(164,671)(391,671){69}
wire w2;    //: /sn:0 {0}(594,314)(846,314)(846,100)(959,100)(959,81){1}
wire w11;    //: /sn:0 {0}(440,201)(411,201)(411,179)(396,179){1}
wire w12;    //: /sn:0 {0}(355,201)(85,201){1}
//: {2}(83,199)(83,134)(195,134)(195,121){3}
//: {4}(83,203)(83,224){5}
//: {6}(85,226)(377,226){7}
//: {8}(83,228)(83,248){9}
//: {10}(85,250)(355,250){11}
//: {12}(83,252)(83,276){13}
//: {14}(85,278)(375,278){15}
//: {16}(83,280)(83,305){17}
//: {18}(85,307)(347,307){19}
//: {20}(83,309)(83,342){21}
//: {22}(85,344)(347,344){23}
//: {24}(83,346)(83,370){25}
//: {26}(85,372)(376,372){27}
//: {28}(83,374)(83,414){29}
//: {30}(85,416)(348,416){31}
//: {32}(83,418)(83,441){33}
//: {34}(85,443)(376,443){35}
//: {36}(83,445)(83,474){37}
//: {38}(85,476)(350,476){39}
//: {40}(83,478)(83,504){41}
//: {42}(85,506)(377,506){43}
//: {44}(83,508)(83,519){45}
//: {46}(85,521)(439,521){47}
//: {48}(83,523)(83,573){49}
//: {50}(85,575)(351,575){51}
//: {52}(83,577)(83,599){53}
//: {54}(85,601)(373,601){55}
//: {56}(83,603)(83,632){57}
//: {58}(85,634)(417,634){59}
//: {60}(83,636)(83,666)(391,666){61}
wire w77;    //: /sn:0 {0}(521,344)(483,344)(483,526)(460,526){1}
wire w13;    //: /sn:0 {0}(368,307)(439,307){1}
wire w27;    //: /sn:0 {0}(594,374)(627,374)(627,158)(694,158)(694,148){1}
//: {2}(696,146)(709,146){3}
//: {4}(713,146)(725,146){5}
//: {6}(729,146)(741,146){7}
//: {8}(745,146)(757,146){9}
//: {10}(761,146)(773,146){11}
//: {12}(777,146)(789,146){13}
//: {14}(793,146)(807,146)(807,143){15}
//: {16}(809,141)(816,141)(816,87)(809,87){17}
//: {18}(807,85)(807,76)(793,76){19}
//: {20}(789,76)(777,76){21}
//: {22}(775,74)(775,77){23}
//: {24}(773,76)(761,76){25}
//: {26}(759,74)(759,65)(758,65)(758,76){27}
//: {28}(757,76)(745,76){29}
//: {30}(741,76)(729,76){31}
//: {32}(727,74)(727,67)(726,67)(726,78){33}
//: {34}(725,76)(713,76){35}
//: {36}(709,76)(695,76)(695,91){37}
//: {38}(711,78)(711,83){39}
//: {40}(743,78)(743,78){41}
//: {42}(791,78)(791,86){43}
//: {44}(807,89)(807,95){45}
//: {46}(807,139)(807,131){47}
//: {48}(791,144)(791,142)(792,142)(792,136){49}
//: {50}(775,148)(775,155)(777,155)(777,145){51}
//: {52}(759,144)(759,156){53}
//: {54}(743,148)(743,165)(742,165)(742,155){55}
//: {56}(727,148)(727,149){57}
//: {58}(711,144)(711,136)(704,136)(704,129){59}
//: {60}(706,127)(711,127){61}
//: {62}(715,127)(727,127){63}
//: {64}(731,127)(743,127){65}
//: {66}(747,127)(759,127){67}
//: {68}(763,127)(775,127){69}
//: {70}(779,127)(791,127){71}
//: {72}(795,127)(808,127)(808,119){73}
//: {74}(793,125)(793,123)(794,123)(794,117){75}
//: {76}(777,129)(777,132)(779,132)(779,122){77}
//: {78}(761,125)(761,127){79}
//: {80}(745,129)(745,137)(746,137)(746,127){81}
//: {82}(729,125)(729,122){83}
//: {84}(713,125)(713,116){85}
//: {86}(702,127)(696,127)(696,112){87}
//: {88}(711,144)(711,139)(711,139)(711,139){89}
//: {90}(694,144)(694,131){91}
wire w33;    //: /sn:0 {0}(369,408)(434,408)(434,327)(439,327){1}
wire w5;    //: /sn:0 {0}(439,526)(390,526)(390,535)(375,535){1}
wire w29;    //: /sn:0 {0}(439,322)(426,322)(426,379)(397,379){1}
wire w9;    //: /sn:0 {0}(397,435)(419,435)(419,457)(438,457){1}
wire w26;    //: /sn:0 {0}(438,467)(413,467)(413,498)(398,498){1}
//: enddecls

  //: joint g165 (w22) @(164, 501) /w:[ 50 49 -1 52 ]
  _GGAND4 #(10) g154 (.I0(w34), .I1(!w30), .I2(!w22), .I3(w12), .Z(w26));   //: @(388,498) /sn:0 /w:[ 9 13 51 43 1 ]
  //: joint g4 (w28) @(734, 370) /w:[ 12 18 11 -1 ]
  //: LED g8 (w28) @(950,157) /sn:0 /w:[ 21 ] /type:0
  //: joint g186 (w22) @(164, 639) /w:[ 66 65 -1 68 ]
  //: joint g140 (w30) @(241, 354) /w:[ 32 34 -1 31 ]
  //: LED g13 (w28) @(885,157) /sn:0 /w:[ 0 ] /type:0
  //: LED g37 (w3) @(1000,190) /sn:0 /w:[ 15 ] /type:0
  //: LED g55 (w27) @(711,132) /sn:0 /w:[ 89 ] /type:0
  //: LED g58 (w27) @(759,149) /sn:0 /w:[ 53 ] /type:0
  //: joint g139 (w22) @(164, 349) /w:[ 30 29 -1 32 ]
  //: joint g112 (w22) @(164, 206) /w:[ 10 9 -1 12 ]
  //: LED g76 (w27) @(775,84) /sn:0 /R:2 /w:[ 23 ] /type:0
  //: joint g111 (w12) @(83, 201) /w:[ 1 2 -1 4 ]
  _GGAND2 #(6) g176 (.I0(w12), .I1(w22), .Z(w24));   //: @(362,578) /sn:0 /w:[ 51 63 1 ]
  //: joint g157 (w30) @(241, 433) /w:[ 20 22 -1 19 ]
  //: joint g163 (w34) @(325, 491) /w:[ 8 10 -1 7 ]
  assign w1 = {w36, w15, w6, w77, w76, w75, w75, w14}; //: CONCAT g1  @(526,339) /sn:0 /w:[ 1 0 0 0 0 0 0 3 0 ] /dr:1 /tp:0 /drp:1
  //: LED g64 (w27) @(807,124) /sn:0 /w:[ 47 ] /type:0
  //: joint g166 (w12) @(83, 506) /w:[ 42 41 -1 44 ]
  //: LED g11 (w28) @(934,157) /sn:0 /w:[ 23 ] /type:0
  //: joint g130 (w22) @(164, 283) /w:[ 22 21 -1 24 ]
  //: joint g121 (w34) @(325, 265) /w:[ 40 42 -1 39 ]
  //: joint g50 (w19) @(917, 142) /w:[ 6 24 5 -1 ]
  //: LED g28 (w3) @(936,190) /sn:0 /w:[ 23 ] /type:0
  //: joint g132 (w34) @(325, 302) /w:[ 36 38 -1 35 ]
  //: LED g19 (w3) @(904,190) /sn:0 /w:[ 27 ] /type:0
  //: joint g113 (w34) @(325, 211) /w:[ 48 50 -1 47 ]
  //: joint g150 (w34) @(325, 387) /w:[ 24 26 -1 23 ]
  //: joint g146 (w30) @(241, 406) /w:[ 24 26 -1 23 ]
  _GGAND2 #(6) g177 (.I0(w12), .I1(w30), .Z(w31));   //: @(384,604) /sn:0 /w:[ 55 5 0 ]
  //: LED g6 (w28) @(966,157) /sn:0 /w:[ 19 ] /type:0
  //: joint g38 (w3) @(703, 415) /w:[ 8 22 7 -1 ]
  //: joint g115 (w22) @(164, 231) /w:[ 14 13 -1 16 ]
  //: joint g53 (w19) @(965, 142) /w:[ 12 18 11 -1 ]
  //: joint g7 (w28) @(750, 370) /w:[ 14 16 13 -1 ]
  //: LED g75 (w27) @(758,83) /sn:0 /R:2 /w:[ 27 ] /type:0
  //: joint g169 (w12) @(83, 521) /w:[ 46 45 -1 48 ]
  //: joint g160 (w34) @(325, 461) /w:[ 12 14 -1 11 ]
  //: joint g135 (w22) @(164, 323) /w:[ 26 25 -1 28 ]
  //: LED g20 (w3) @(968,190) /sn:0 /w:[ 19 ] /type:0
  //: LED g31 (w3) @(920,190) /sn:0 /w:[ 25 ] /type:0
  _GGOR6 #(14) g149 (.I0(w8), .I1(w13), .I2(w21), .I3(w25), .I4(w29), .I5(w33), .Z(w75));   //: @(450,314) /sn:0 /w:[ 1 1 1 0 0 1 5 ]
  _GGAND3 #(8) g124 (.I0(w34), .I1(w12), .I2(!w30), .Z(w13));   //: @(358,307) /sn:0 /w:[ 37 19 41 0 ]
  //: LED g39 (w19) @(901,120) /sn:0 /w:[ 27 ] /type:0
  //: joint g68 (w27) @(727, 76) /w:[ 31 32 34 -1 ]
  //: joint g48 (w19) @(981, 142) /w:[ 14 16 13 -1 ]
  //: joint g17 (w3) @(687, 415) /w:[ 6 24 5 -1 ]
  //: joint g25 (w3) @(719, 415) /w:[ 10 20 9 -1 ]
  //: joint g179 (w12) @(83, 575) /w:[ 50 49 -1 52 ]
  //: joint g52 (w19) @(949, 142) /w:[ 10 20 9 -1 ]
  //: joint g106 (w34) @(325, 150) /w:[ 56 58 -1 55 ]
  //: joint g107 (w22) @(164, 155) /w:[ 1 2 -1 4 ]
  //: joint g174 (w34) @(325, 537) /w:[ 4 6 -1 3 ]
  //: joint g83 (w27) @(745, 127) /w:[ 66 -1 65 80 ]
  //: joint g100 (w27) @(694, 146) /w:[ 2 90 -1 1 ]
  //: LED g14 (w28) @(998,157) /sn:0 /w:[ 15 ] /type:0
  //: DIP g193 (w0) @(209,77) /sn:0 /w:[ 1 ] /st:11 /dn:1
  //: LED g44 (w19) @(981,120) /sn:0 /w:[ 17 ] /type:0
  //: joint g47 (w27) @(727, 146) /w:[ 6 -1 5 56 ]
  //: LED g80 (w27) @(746,120) /sn:0 /w:[ 81 ] /type:0
  //: joint g94 (w27) @(704, 127) /w:[ 60 -1 86 59 ]
  //: joint g172 (w22) @(164, 532) /w:[ 54 53 -1 56 ]
  //: joint g159 (w12) @(83, 443) /w:[ 34 33 -1 36 ]
  //: joint g21 (w3) @(751, 415) /w:[ 14 16 13 -1 ]
  //: joint g84 (w27) @(761, 127) /w:[ 68 78 67 -1 ]
  _GGAND4 #(10) g105 (.I0(w12), .I1(!w22), .I2(!w30), .I3(!w34), .Z(w23));   //: @(366,257) /sn:0 /w:[ 11 19 49 41 1 ]
  //: joint g155 (w12) @(83, 476) /w:[ 38 37 -1 40 ]
  //: joint g141 (w34) @(325, 359) /w:[ 28 30 -1 27 ]
  assign {w27, w3, w28, w19, w32, w4, w2, w35} = w1; //: CONCAT g23  @(589,339) /sn:0 /R:2 /w:[ 0 29 29 29 1 0 0 0 0 ] /dr:0 /tp:0 /drp:0
  //: LED g41 (w19) @(933,120) /sn:0 /w:[ 23 ] /type:0
  //: joint g151 (w75) @(491, 314) /w:[ 2 -1 4 1 ]
  //: LED g40 (w19) @(917,120) /sn:0 /w:[ 25 ] /type:0
  //: joint g54 (w27) @(775, 146) /w:[ 12 -1 11 50 ]
  //: joint g93 (w27) @(713, 127) /w:[ 62 84 61 -1 ]
  //: joint g116 (w30) @(241, 236) /w:[ 52 54 -1 51 ]
  _GGAND3 #(8) g123 (.I0(!w12), .I1(!w22), .I2(w30), .Z(w8));   //: @(386,283) /sn:0 /w:[ 15 23 45 0 ]
  _GGOR3 #(8) g167 (.I0(w9), .I1(w18), .I2(w26), .Z(w76));   //: @(449,462) /sn:0 /w:[ 1 0 0 1 ]
  //: LED g0 (w4) @(902,74) /sn:0 /w:[ 1 ] /type:0
  //: LED g26 (w3) @(984,190) /sn:0 /w:[ 17 ] /type:0
  //: joint g46 (w27) @(711, 146) /w:[ 4 58 3 88 ]
  //: joint g90 (w27) @(729, 127) /w:[ 64 82 63 -1 ]
  //: LED g82 (w27) @(761,120) /sn:0 /w:[ 79 ] /type:0
  //: joint g136 (w30) @(241, 328) /w:[ 36 38 -1 35 ]
  _GGAND4 #(10) g128 (.I0(!w34), .I1(w30), .I2(w22), .I3(w12), .Z(w33));   //: @(359,408) /sn:0 /w:[ 21 25 39 31 0 ]
  //: joint g173 (w22) @(164, 554) /w:[ 58 57 -1 60 ]
  //: LED g33 (w32) @(985,74) /sn:0 /w:[ 0 ] /type:0
  //: joint g91 (w27) @(777, 127) /w:[ 70 -1 69 76 ]
  //: joint g49 (w19) @(933, 142) /w:[ 8 22 7 -1 ]
  //: joint g137 (w34) @(325, 333) /w:[ 32 34 -1 31 ]
  //: LED g61 (w27) @(742,148) /sn:0 /w:[ 55 ] /type:0
  //: joint g158 (w22) @(164, 438) /w:[ 42 41 -1 44 ]
  //: joint g51 (w19) @(901, 142) /w:[ 4 26 3 -1 ]
  //: joint g3 (w28) @(686, 370) /w:[ 6 24 5 -1 ]
  //: joint g86 (w27) @(793, 127) /w:[ 72 74 71 -1 ]
  //: LED g89 (w27) @(779,115) /sn:0 /w:[ 77 ] /type:0
  //: joint g2 (w28) @(670, 370) /w:[ 4 26 3 -1 ]
  //: joint g65 (w27) @(743, 146) /w:[ 8 -1 7 54 ]
  //: LED g77 (w27) @(807,102) /sn:0 /R:2 /w:[ 45 ] /type:0
  //: joint g110 (w34) @(325, 184) /w:[ 52 54 -1 51 ]
  //: joint g156 (w34) @(325, 428) /w:[ 16 18 -1 15 ]
  //: joint g148 (w12) @(83, 416) /w:[ 30 29 -1 32 ]
  //: joint g147 (w22) @(164, 411) /w:[ 38 37 -1 40 ]
  //: joint g59 (w27) @(759, 146) /w:[ 10 52 9 -1 ]
  _GGAND4 #(10) g153 (.I0(!w34), .I1(w30), .I2(w22), .I3(w12), .Z(w18));   //: @(361,468) /sn:0 /w:[ 13 17 47 39 1 ]
  //: LED g72 (w27) @(743,85) /sn:0 /R:2 /w:[ 41 ] /type:0
  //: joint g99 (w3) @(654, 415) /w:[ 2 1 28 -1 ]
  //: joint g98 (w28) @(653, 370) /w:[ 2 1 28 -1 ]
  //: joint g182 (w30) @(241, 606) /w:[ 4 6 -1 3 ]
  //: joint g161 (w30) @(241, 466) /w:[ 16 18 -1 15 ]
  //: joint g16 (w3) @(671, 415) /w:[ 4 26 3 -1 ]
  //: joint g96 (w27) @(807, 141) /w:[ 16 46 -1 15 ]
  _GGAND4 #(10) g183 (.I0(w12), .I1(w22), .I2(w30), .I3(w34), .Z(w15));   //: @(428,641) /sn:0 /w:[ 59 67 0 0 1 ]
  _GGAND4 #(10) g152 (.I0(!w34), .I1(!w30), .I2(w22), .I3(!w12), .Z(w9));   //: @(387,435) /sn:0 /w:[ 17 21 43 35 0 ]
  _GGAND3 #(8) g103 (.I0(!w12), .I1(w22), .I2(!w34), .Z(w16));   //: @(366,206) /sn:0 /w:[ 0 11 49 1 ]
  _GGOR5 #(12) g122 (.I0(w7), .I1(w11), .I2(w16), .I3(w20), .I4(w23), .Z(w14));   //: @(451,206) /sn:0 /w:[ 1 0 0 0 0 1 ]
  //: LED g10 (w28) @(982,157) /sn:0 /w:[ 17 ] /type:0
  //: LED g78 (w27) @(695,98) /sn:0 /R:2 /w:[ 37 ] /type:0
  //: LED g87 (w27) @(729,115) /sn:0 /w:[ 83 ] /type:0
  _GGAND2 #(6) g171 (.I0(w22), .I1(w30), .Z(w17));   //: @(392,557) /sn:0 /w:[ 59 9 1 ]
  //: joint g129 (w12) @(83, 278) /w:[ 14 13 -1 16 ]
  //: LED g32 (w35) @(932,74) /sn:0 /w:[ 1 ] /type:0
  //: joint g187 (w30) @(241, 644) /w:[ 1 2 -1 60 ]
  _GGAND3 #(8) g102 (.I0(w22), .I1(w30), .I2(!w34), .Z(w11));   //: @(386,179) /sn:0 /w:[ 7 57 53 1 ]
  //: LED g69 (w27) @(791,93) /sn:0 /R:2 /w:[ 43 ] /type:0
  //: joint g143 (w22) @(164, 377) /w:[ 34 33 -1 36 ]
  //: joint g9 (w28) @(718, 370) /w:[ 10 20 9 -1 ]
  //: joint g57 (w27) @(791, 146) /w:[ 14 48 13 -1 ]
  //: joint g119 (w22) @(164, 255) /w:[ 18 17 -1 20 ]
  //: joint g71 (w27) @(711, 76) /w:[ 35 -1 36 38 ]
  //: joint g15 (w28) @(702, 370) /w:[ 8 22 7 -1 ]
  //: joint g142 (w12) @(83, 372) /w:[ 26 25 -1 28 ]
  //: joint g162 (w22) @(164, 471) /w:[ 46 45 -1 48 ]
  _GGAND4 #(10) g127 (.I0(w12), .I1(!w22), .I2(!w30), .I3(!w34), .Z(w29));   //: @(387,379) /sn:0 /w:[ 27 35 29 25 1 ]
  //: joint g67 (w27) @(775, 76) /w:[ 21 22 24 -1 ]
  //: joint g131 (w30) @(241, 288) /w:[ 44 46 -1 43 ]
  //: LED g43 (w19) @(965,120) /sn:0 /w:[ 19 ] /type:0
  //: LED g62 (w27) @(727,142) /sn:0 /w:[ 57 ] /type:0
  //: joint g145 (w34) @(325, 401) /w:[ 20 22 -1 19 ]
  //: joint g73 (w27) @(743, 76) /w:[ 30 40 29 -1 ]
  //: LED g88 (w27) @(696,105) /sn:0 /w:[ 87 ] /type:0
  _GGAND4 #(10) g104 (.I0(w12), .I1(w22), .I2(!w30), .I3(w34), .Z(w20));   //: @(388,233) /sn:0 /w:[ 7 15 53 45 1 ]
  //: joint g138 (w12) @(83, 344) /w:[ 22 21 -1 24 ]
  //: LED g42 (w19) @(949,120) /sn:0 /w:[ 21 ] /type:0
  //: LED g63 (w27) @(694,124) /sn:0 /w:[ 91 ] /type:0
  //: joint g180 (w12) @(83, 601) /w:[ 54 53 -1 56 ]
  //: joint g188 (w34) @(325, 649) /w:[ 1 2 -1 60 ]
  //: LED g74 (w27) @(711,90) /sn:0 /R:2 /w:[ 39 ] /type:0
  //: joint g109 (w30) @(241, 179) /w:[ 56 58 -1 55 ]
  //: joint g175 (w30) @(241, 559) /w:[ 8 10 -1 7 ]
  //: joint g133 (w12) @(83, 307) /w:[ 18 17 -1 20 ]
  //: LED g5 (w28) @(902,157) /sn:0 /w:[ 27 ] /type:0
  //: LED g56 (w27) @(777,138) /sn:0 /w:[ 51 ] /type:0
  _GGOR3 #(8) g168 (.I0(w12), .I1(w5), .I2(w17), .Z(w77));   //: @(450,526) /sn:0 /w:[ 47 0 0 1 ]
  //: joint g181 (w22) @(164, 580) /w:[ 62 61 -1 64 ]
  //: joint g79 (w27) @(759, 76) /w:[ 25 26 28 -1 ]
  //: joint g95 (w27) @(807, 87) /w:[ 17 18 -1 44 ]
  //: joint g117 (w34) @(325, 241) /w:[ 44 46 -1 43 ]
  assign {w12, w22, w30, w34} = w0; //: CONCAT g194  @(210,116) /sn:0 /R:1 /w:[ 3 3 59 59 0 ] /dr:0 /tp:0 /drp:0
  //: LED g92 (w27) @(794,110) /sn:0 /w:[ 75 ] /type:0
  //: LED g85 (w27) @(808,112) /sn:0 /w:[ 73 ] /type:0
  //: LED g24 (w2) @(959,74) /sn:0 /w:[ 1 ] /type:0
  //: LED g36 (w3) @(887,190) /sn:0 /w:[ 0 ] /type:0
  _GGAND3 #(8) g125 (.I0(w22), .I1(!w30), .I2(!w34), .Z(w21));   //: @(387,328) /sn:0 /w:[ 27 37 33 0 ]
  //: joint g144 (w30) @(241, 382) /w:[ 28 30 -1 27 ]
  _GGOR2 #(6) g178 (.I0(w24), .I1(w31), .Z(w6));   //: @(453,596) /sn:0 /w:[ 0 1 1 ]
  _GGAND2 #(6) g101 (.I0(w34), .I1(!w22), .Z(w7));   //: @(364,153) /sn:0 /w:[ 57 0 0 ]
  //: LED g81 (w27) @(713,109) /sn:0 /w:[ 85 ] /type:0
  //: LED g60 (w27) @(792,129) /sn:0 /w:[ 49 ] /type:0
  _GGAND4 #(10) g126 (.I0(!w12), .I1(w22), .I2(w30), .I3(w34), .Z(w25));   //: @(358,351) /sn:0 /w:[ 23 31 33 29 1 ]
  //: LED g70 (w27) @(726,85) /sn:0 /R:2 /w:[ 33 ] /type:0
  //: LED g22 (w3) @(952,190) /sn:0 /w:[ 21 ] /type:0
  //: LED g45 (w19) @(997,120) /sn:0 /w:[ 15 ] /type:0
  //: LED g35 (w19) @(884,120) /sn:0 /w:[ 0 ] /type:0
  _GGAND2 #(6) g170 (.I0(w22), .I1(w34), .Z(w5));   //: @(365,535) /sn:0 /w:[ 55 5 1 ]
  //: joint g185 (w12) @(83, 634) /w:[ 58 57 -1 60 ]
  //: joint g120 (w30) @(241, 260) /w:[ 48 50 -1 47 ]
  //: joint g114 (w12) @(83, 226) /w:[ 6 5 -1 8 ]
  //: joint g66 (w27) @(791, 76) /w:[ 19 -1 20 42 ]
  //: joint g97 (w19) @(884, 142) /w:[ 2 1 -1 28 ]
  _GGAND4 #(8) g184 (.I0(!w12), .I1(!w22), .I2(!w30), .I3(!w34), .Z(w36));   //: @(402,673) /sn:0 /w:[ 61 69 61 61 1 ]
  //: joint g18 (w3) @(735, 415) /w:[ 12 18 11 -1 ]
  //: LED g12 (w28) @(918,157) /sn:0 /w:[ 25 ] /type:0
  //: joint g164 (w30) @(241, 496) /w:[ 12 14 -1 11 ]
  //: joint g108 (w22) @(164, 174) /w:[ 6 5 -1 8 ]
  //: joint g118 (w12) @(83, 250) /w:[ 10 9 -1 12 ]
  //: joint g134 (w30) @(241, 312) /w:[ 40 42 -1 39 ]

endmodule
//: /netlistEnd

