//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
input Clock;    //: /sn:0 {0}(123,435)(273,435){1}
//: {2}(277,435)(366,435){3}
//: {4}(370,435)(551,435)(551,324){5}
//: {6}(368,433)(368,324){7}
//: {8}(275,433)(275,324){9}
input [3:0] Din;    //: /sn:0 {0}(#:109,338)(#:177,338){1}
input Enable;    //: {0}(189,219)(164,219)(164,216)(52:141,216){1}
output [3:0] Dout;    //: /sn:0 {0}(#:663,314)(705,314){1}
input Reset;    //: /sn:0 {0}(189,176)(155,176)(155,177)(140,177){1}
wire w6;    //: /sn:0 {0}(657,329)(610,329)(610,235)(295,235)(295,303)(291,303){1}
wire w7;    //: /sn:0 {0}(445,307)(427,307)(427,343)(183,343){1}
wire w14;    //: /sn:0 {0}(384,303)(396,303)(396,247)(632,247)(632,319)(657,319){1}
wire w15;    //: /sn:0 {0}(384,313)(399,313){1}
wire w4;    //: /sn:0 {0}(259,308)(198,308)(198,323)(183,323){1}
wire w3;    //: /sn:0 {0}(205,219)(278,219){1}
//: {2}(282,219)(371,219){3}
//: {4}(375,219)(464,219){5}
//: {6}(468,219)(556,219)(556,292){7}
//: {8}(466,221)(466,291){9}
//: {10}(373,221)(373,292){11}
//: {12}(280,221)(280,292){13}
wire w21;    //: /sn:0 {0}(477,312)(492,312){1}
wire w20;    //: /sn:0 {0}(477,302)(487,302)(487,261)(624,261)(624,309)(657,309){1}
wire w1;    //: /sn:0 {0}(205,176)(361,176){1}
//: {2}(365,176)(454,176){3}
//: {4}(458,176)(546,176)(546,292){5}
//: {6}(456,178)(456,291){7}
//: {8}(363,178)(363,292){9}
wire w25;    //: /sn:0 {0}(461,436)(461,323){1}
wire w8;    //: /sn:0 {0}(535,308)(512,308)(512,353)(183,353){1}
wire w12;    //: /sn:0 {0}(270,179)(270,292){1}
wire w27;    //: /sn:0 {0}(567,313)(582,313){1}
wire w5;    //: /sn:0 {0}(352,308)(332,308)(332,333)(183,333){1}
wire w9;    //: /sn:0 {0}(291,313)(306,313){1}
wire w26;    //: /sn:0 {0}(567,303)(642,303)(642,299)(657,299){1}
//: enddecls

  _GGFF #(10, 10, 20) g8 (.Q(w14), ._Q(w15), .D(w5), .EN(w3), .CLR(w1), .CK(Clock));   //: @(368,308) /sn:0 /w:[ 0 0 0 11 9 7 ] /mi:0
  //: IN g4 (Din) @(107,338) /sn:0 /w:[ 0 ]
  //: joint g13 (w3) @(280, 219) /w:[ 2 -1 1 12 ]
  _GGNBUF #(2) g3 (.I(Enable), .Z(w3));   //: @(195,219) /sn:0 /w:[ 0 0 ]
  _GGNBUF #(2) g2 (.I(Reset), .Z(w1));   //: @(195,176) /sn:0 /w:[ 0 0 ]
  //: IN g1 (Enable) @(139,216) /sn:0 /w:[ 1 ]
  //: joint g16 (Clock) @(368, 435) /w:[ 4 6 3 -1 ]
  //: joint g11 (w1) @(456, 176) /w:[ 4 -1 3 6 ]
  _GGFF #(10, 10, 20) g10 (.Q(w26), ._Q(w27), .D(w8), .EN(w3), .CLR(w1), .CK(Clock));   //: @(551,308) /sn:0 /w:[ 0 0 0 7 5 5 ] /mi:0
  //: OUT g19 (Dout) @(702,314) /sn:0 /w:[ 1 ]
  assign {w8, w7, w5, w4} = Din; //: CONCAT g6  @(178,338) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  _GGFF #(10, 10, 20) g9 (.Q(w20), ._Q(w21), .D(w7), .EN(w3), .CLR(w1), .CK(w25));   //: @(461,307) /sn:0 /w:[ 0 0 0 9 7 1 ] /mi:0
  _GGFF #(10, 10, 20) g7 (.Q(w6), ._Q(w9), .D(w4), .EN(w3), .CLR(w12), .CK(Clock));   //: @(275,308) /sn:0 /w:[ 1 0 0 13 1 9 ] /mi:0
  //: joint g15 (w3) @(466, 219) /w:[ 6 -1 5 8 ]
  //: joint g17 (Clock) @(275, 435) /w:[ 2 8 1 -1 ]
  //: joint g14 (w3) @(373, 219) /w:[ 4 -1 3 10 ]
  //: IN g5 (Clock) @(121,435) /sn:0 /w:[ 0 ]
  //: IN g0 (Reset) @(138,177) /sn:0 /w:[ 1 ]
  assign Dout = {w26, w20, w14, w6}; //: CONCAT g18  @(662,314) /sn:0 /w:[ 0 1 1 1 0 ] /dr:0 /tp:0 /drp:1
  //: joint g12 (w1) @(363, 176) /w:[ 2 -1 1 8 ]

endmodule
//: /netlistEnd

