//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "ALU_8functions.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [7:0] B;    //: /sn:0 {0}(#:200,350)(200,257){1}
//: {2}(202,255)(#:212,255)(212,264)(341,264){3}
//: {4}(200,253)(200,237){5}
//: {6}(202,235)(#:212,235)(212,239)(338,239){7}
//: {8}(200,233)(200,188){9}
//: {10}(202,186)(335,186){11}
//: {12}(200,184)(200,170){13}
//: {14}(202,168)(#:229,168)(229,276)(324,276)(324,292)(341,292){15}
//: {16}(200,166)(200,154){17}
//: {18}(202,152)(338,152){19}
//: {20}(200,150)(200,101)(247,101)(#:247,69){21}
reg [7:0] A;    //: /sn:0 {0}(#:120,68)(120,119){1}
//: {2}(122,121)(419,121)(419,135)(496,135)(496,176)(534,176){3}
//: {4}(120,123)(120,156){5}
//: {6}(122,158)(#:132,158)(132,157)(338,157){7}
//: {8}(120,160)(120,187){9}
//: {10}(122,189)(#:132,189)(132,191)(335,191){11}
//: {12}(120,191)(120,214){13}
//: {14}(122,216)(340,216){15}
//: {16}(120,218)(120,245){17}
//: {18}(122,247)(#:132,247)(132,244)(338,244){19}
//: {20}(120,249)(120,267){21}
//: {22}(122,269)(341,269){23}
//: {24}(120,271)(120,280)(148,280){25}
//: {26}(152,280)(216,280)(216,350){27}
//: {28}(#:150,282)(150,297)(341,297){29}
reg w21;    //: /sn:0 {0}(534,144)(482,144)(482,44)(460,44){1}
reg w23;    //: /sn:0 {0}(521,43)(531,43)(531,58)(519,58)(519,160)(534,160){1}
reg w22;    //: /sn:0 {0}(397,43)(407,43)(407,58)(384,58)(384,87)(471,87)(471,128)(534,128){1}
wire [7:0] w6;    //: /sn:0 {0}(#:356,189)(428,189)(428,256)(534,256){1}
wire [7:0] w7;    //: /sn:0 {0}(#:362,295)(453,295)(453,272)(534,272){1}
wire [7:0] w14;    //: /sn:0 {0}(#:362,267)(500,267)(500,208)(534,208){1}
wire [7:0] w4;    //: /sn:0 {0}(#:356,216)(519,216)(519,240)(534,240){1}
wire [7:0] w0;    //: /sn:0 {0}(#:699,103)(699,128)(596,128){1}
wire [7:0] w1;    //: /sn:0 {0}(#:216,450)(216,553)(291,553)(291,381)(420,381)(420,288)(534,288){1}
wire [7:0] w8;    //: /sn:0 {0}(#:359,242)(484,242)(484,192)(534,192){1}
wire [7:0] w2;    //: /sn:0 {0}(200,450)(200,507)(#:104,507)(104,441){1}
wire [7:0] w13;    //: /sn:0 {0}(#:359,155)(442,155)(442,224)(534,224){1}
//: enddecls

  //: joint g4 (A) @(120, 121) /w:[ 2 1 -1 4 ]
  _GGOR2x8 #(6) g8 (.I0(B), .I1(A), .Z(w6));   //: @(346,189) /sn:0 /w:[ 11 11 0 ]
  //: LED g3 (w0) @(699,96) /sn:0 /w:[ 0 ] /type:3
  //: comment g13 @(271,136) /sn:0
  //: /line:"A AND B"
  //: /line:""
  //: /end
  //: comment g34 @(252,222) /sn:0
  //: /line:"1-"
  //: /end
  //: comment g37 @(226,472) /sn:0
  //: /line:"7-"
  //: /end
  //: DIP g2 (B) @(247,59) /sn:0 /w:[ 21 ] /st:0 /dn:1
  //: LED g1 (w2) @(104,434) /sn:0 /w:[ 1 ] /type:0
  //: DIP A (A) @(120,58) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGNBUF8 #(2) g11 (.I(A), .Z(w4));   //: @(346,216) /sn:0 /w:[ 15 0 ]
  _GGXOR2x8 #(8) g16 (.I0(B), .I1(A), .Z(w8));   //: @(349,242) /sn:0 /w:[ 7 19 0 ]
  //: joint g10 (A) @(120, 189) /w:[ 10 9 -1 12 ]
  //: comment g28 @(266,281) /sn:0
  //: /line:"A NOR B"
  //: /end
  //: comment g19 @(267,226) /sn:0
  //: /line:"A XOR B"
  //: /end
  //: joint g27 (A) @(150, 280) /w:[ 26 -1 25 28 ]
  //: comment g32 @(254,135) /sn:0
  //: /line:"3-"
  //: /end
  //: joint g6 (B) @(200, 152) /w:[ 18 20 -1 17 ]
  mux g38 (.s0(w22), .s1(w21), .s2(w23), .x0(A), .x1(w8), .x2(w14), .x3(w13), .x4(w4), .x5(w6), .x6(w7), .x7(w1), .y0(w0));   //: @(535, 112) /sz:(60, 192) /sn:0 /p:[ Li0>1 Li1>0 Li2>1 Li3>3 Li4>1 Li5>1 Li6>1 Li7>1 Li8>1 Li9>1 Li10>1 Ro0<1 ]
  //: joint g7 (A) @(120, 158) /w:[ 6 5 -1 8 ]
  //: joint g9 (B) @(200, 186) /w:[ 10 12 -1 9 ]
  //: comment g15 @(275,204) /sn:0
  //: /line:"NOT A"
  //: /end
  _GGNAND2x8 #(4) g20 (.I0(B), .I1(A), .Z(w14));   //: @(352,267) /sn:0 /w:[ 3 23 0 ]
  //: comment g31 @(258,170) /sn:0
  //: /line:"5-"
  //: /end
  //: SWITCH g39 (w21) @(443,44) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: joint g17 (B) @(200, 235) /w:[ 6 8 -1 5 ]
  _GGNOR2x8 #(4) g25 (.I0(B), .I1(A), .Z(w7));   //: @(352,295) /sn:0 /w:[ 15 29 0 ]
  //: comment g29 @(244,473) /sn:0
  //: /line:"A + B"
  //: /end
  _GGAND2x8 #(6) g5 (.I0(B), .I1(A), .Z(w13));   //: @(349,155) /sn:0 /w:[ 19 7 0 ]
  //: comment g14 @(272,174) /sn:0
  //: /line:"A OR B"
  //: /end
  //: joint g21 (B) @(200, 255) /w:[ 2 4 -1 1 ]
  //: comment g24 @(284,106) /sn:0
  //: /line:"A"
  //: /end
  //: comment g36 @(246,279) /sn:0
  //: /line:"6-"
  //: /end
  //: comment g23 @(264,251) /sn:0
  //: /line:"A NAND B"
  //: /end
  //: SWITCH g41 (w23) @(504,43) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g40 (w22) @(380,43) /sn:0 /w:[ 0 ] /st:0 /dn:1
  adder g0 (.a0(A), .b0(B), .res(w1), .sign(w2));   //: @(184, 351) /sz:(48, 98) /R:3 /sn:0 /p:[ Ti0>27 Ti1>0 Bo0<0 Bo1<0 ]
  //: joint g22 (A) @(120, 269) /w:[ 22 21 -1 24 ]
  //: joint g26 (B) @(200, 168) /w:[ 14 16 -1 13 ]
  //: comment g35 @(248,250) /sn:0
  //: /line:"2-"
  //: /end
  //: joint g12 (A) @(120, 216) /w:[ 14 13 -1 16 ]
  //: joint g18 (A) @(120, 247) /w:[ 18 17 -1 20 ]
  //: comment g30 @(267,105) /sn:0
  //: /line:"0-"
  //: /end
  //: comment g33 @(257,200) /sn:0
  //: /line:"4-"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin mux
module mux(x4, x3, x2, x1, s1, x6, x7, s2, y0, x5, x0, s0);
//: interface  /sz:(60, 192) /bd:[ Li0>s0(16/192) Li1>s1(32/192) Li2>s2(48/192) Li3>x0[7:0](64/192) Li4>x1[7:0](80/192) Li5>x2[7:0](96/192) Li6>x3[7:0](112/192) Li7>x4[7:0](128/192) Li8>x5[7:0](144/192) Li9>x6[7:0](160/192) Li10>x7[7:0](176/192) Ro0<y0[7:0](16/192) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [7:0] x1;    //: /sn:0 {0}(#:63,115)(364,115)(364,113)(397,113){1}
input s2;    //: /sn:0 {0}(396,298)(279,298){1}
//: {2}(277,296)(277,257){3}
//: {4}(279,255)(396,255){5}
//: {6}(277,253)(277,217){7}
//: {8}(279,215)(339,215){9}
//: {10}(277,213)(277,181){11}
//: {12}(279,179)(289,179)(289,182)(307,182){13}
//: {14}(277,177)(277,146){15}
//: {16}(279,144)(309,144){17}
//: {18}(277,142)(277,81)(301,81){19}
//: {20}(277,300)(277,343){21}
//: {22}(279,345)(289,345)(289,338)(396,338){23}
//: {24}(277,347)(277,385){25}
//: {26}(279,387)(289,387)(289,382)(396,382){27}
//: {28}(277,389)(277,488)(271,488){29}
input s0;    //: /sn:0 {0}(193,431)(204,431)(204,374){1}
//: {2}(206,372)(396,372){3}
//: {4}(204,370)(204,338){5}
//: {6}(206,336)(216,336)(216,327)(309,327){7}
//: {8}(204,334)(204,290){9}
//: {10}(206,288)(396,288){11}
//: {12}(204,286)(204,247){13}
//: {14}(206,245)(216,245)(216,240)(302,240){15}
//: {16}(204,243)(204,208){17}
//: {18}(206,206)(216,206)(216,205)(397,205){19}
//: {20}(204,204)(204,169){21}
//: {22}(206,167)(216,167)(216,163)(310,163){23}
//: {24}(204,165)(204,126){25}
//: {26}(206,124)(216,124)(216,118)(397,118){27}
//: {28}(204,122)(204,49)(300,49){29}
input [7:0] x0;    //: /sn:0 {0}(#:63,78)(322,78)(322,71)(396,71){1}
output [7:0] y0;    //: /sn:0 {0}(658,222)(#:601,222){1}
input [7:0] x7;    //: /sn:0 {0}(#:70,338)(132,338)(132,367)(396,367){1}
input s1;    //: /sn:0 {0}(396,333)(255,333)(255,337)(245,337){1}
//: {2}(243,335)(243,295){3}
//: {4}(245,293)(255,293)(255,294)(296,294){5}
//: {6}(243,291)(243,254){7}
//: {8}(245,252)(255,252)(255,250)(303,250){9}
//: {10}(243,250)(243,213){11}
//: {12}(245,211)(255,211)(255,210)(397,210){13}
//: {14}(243,209)(243,170){15}
//: {16}(245,168)(255,168)(255,167)(398,167){17}
//: {18}(243,166)(243,130){19}
//: {20}(245,128)(308,128){21}
//: {22}(243,126)(243,65)(301,65){23}
//: {24}(243,339)(243,379){25}
//: {26}(245,381)(255,381)(255,377)(396,377){27}
//: {28}(243,383)(243,461)(224,461){29}
input [7:0] x4;    //: /sn:0 {0}(#:67,228)(385,228)(385,240)(396,240){1}
input [7:0] x6;    //: /sn:0 {0}(#:70,302)(179,302)(179,323)(396,323){1}
input [7:0] x3;    //: /sn:0 {0}(#:67,191)(386,191)(386,200)(397,200){1}
input [7:0] x5;    //: /sn:0 {0}(#:68,263)(308,263)(308,283)(396,283){1}
input [7:0] x2;    //: /sn:0 {0}(#:65,152)(387,152)(387,157)(398,157){1}
wire w7;    //: /sn:0 {0}(324,128)(374,128)(374,123)(397,123){1}
wire [7:0] w14;    //: /sn:0 {0}(#:419,164)(522,164)(522,215)(#:580,215){1}
wire w4;    //: /sn:0 {0}(317,81)(339,81)(339,86)(396,86){1}
wire [7:0] w19;    //: /sn:0 {0}(#:418,207)(480,207)(480,220)(#:580,220){1}
wire w3;    //: /sn:0 {0}(317,65)(354,65)(354,81)(396,81){1}
wire w37;    //: /sn:0 {0}(319,250)(396,250){1}
wire [7:0] w34;    //: /sn:0 {0}(#:417,330)(522,330)(522,235)(#:580,235){1}
wire w31;    //: /sn:0 {0}(325,327)(377,327)(377,328)(396,328){1}
wire [7:0] w24;    //: /sn:0 {0}(#:417,290)(514,290)(514,230)(#:580,230){1}
wire w36;    //: /sn:0 {0}(318,240)(381,240)(381,245)(396,245){1}
wire w1;    //: /sn:0 {0}(316,49)(381,49)(381,76)(396,76){1}
wire w8;    //: /sn:0 {0}(325,144)(382,144)(382,128)(397,128){1}
wire w18;    //: /sn:0 {0}(355,215)(397,215){1}
wire w22;    //: /sn:0 {0}(312,294)(368,294)(368,293)(396,293){1}
wire [7:0] w2;    //: /sn:0 {0}(#:417,78)(565,78)(565,205)(580,205){1}
wire w11;    //: /sn:0 {0}(326,163)(383,163)(383,162)(398,162){1}
wire w13;    //: /sn:0 {0}(323,182)(383,182)(383,172)(398,172){1}
wire [7:0] w29;    //: /sn:0 {0}(#:417,374)(533,374)(533,240)(#:580,240){1}
wire [7:0] w9;    //: /sn:0 {0}(#:418,120)(543,120)(543,210)(580,210){1}
wire [7:0] w39;    //: /sn:0 {0}(#:417,247)(509,247)(509,225)(#:580,225){1}
//: enddecls

  //: IN g4 (x4) @(65,228) /sn:0 /w:[ 0 ]
  _GGAND4x8 #(10) g8 (.I0(x0), .I1({8{w1}}), .I2({8{w3}}), .I3({8{w4}}), .Z(w2));   //: @(407,78) /sn:0 /w:[ 1 1 1 1 0 ]
  //: IN g3 (x3) @(65,191) /sn:0 /w:[ 0 ]
  _GGAND4x8 #(10) g13 (.I0(x7), .I1({8{s0}}), .I2({8{s1}}), .I3({8{s2}}), .Z(w29));   //: @(407,374) /sn:0 /w:[ 1 3 27 27 0 ]
  //: joint g34 (s1) @(243, 168) /w:[ 16 18 -1 15 ]
  _GGNBUF #(2) g37 (.I(s2), .Z(w18));   //: @(345,215) /sn:0 /w:[ 9 0 ]
  //: joint g51 (s2) @(277, 298) /w:[ 1 2 -1 20 ]
  //: IN g2 (x2) @(63,152) /sn:0 /w:[ 0 ]
  //: IN g1 (x1) @(61,115) /sn:0 /w:[ 0 ]
  _GGAND4x8 #(10) g11 (.I0(x3), .I1({8{s0}}), .I2({8{s1}}), .I3({8{w18}}), .Z(w19));   //: @(408,207) /sn:0 /w:[ 1 19 13 1 0 ]
  _GGOR8x8 #(18) g16 (.I0(w2), .I1(w9), .I2(w14), .I3(w19), .I4(w39), .I5(w24), .I6(w34), .I7(w29), .Z(y0));   //: @(591,222) /sn:0 /w:[ 1 1 1 1 1 1 1 1 1 ]
  _GGAND4x8 #(10) g10 (.I0(x2), .I1({8{w11}}), .I2({8{s1}}), .I3({8{w13}}), .Z(w14));   //: @(409,164) /sn:0 /w:[ 1 1 17 1 0 ]
  _GGNBUF #(2) g28 (.I(s2), .Z(w8));   //: @(315,144) /sn:0 /w:[ 17 0 ]
  _GGNBUF #(2) g50 (.I(s1), .Z(w22));   //: @(302,294) /sn:0 /w:[ 5 0 ]
  //: IN g19 (s1) @(222,461) /sn:0 /w:[ 29 ]
  _GGNBUF #(2) g27 (.I(s1), .Z(w7));   //: @(314,128) /sn:0 /w:[ 21 0 ]
  _GGNBUF #(2) g32 (.I(s0), .Z(w11));   //: @(316,163) /sn:0 /w:[ 23 0 ]
  //: IN g6 (x6) @(68,302) /sn:0 /w:[ 0 ]
  //: joint g38 (s2) @(277, 215) /w:[ 8 10 -1 7 ]
  //: IN g7 (x7) @(68,338) /sn:0 /w:[ 0 ]
  _GGAND4x8 #(10) g9 (.I0(x1), .I1({8{s0}}), .I2({8{w7}}), .I3({8{w8}}), .Z(w9));   //: @(408,120) /sn:0 /w:[ 1 27 1 1 0 ]
  //: joint g53 (s0) @(204, 288) /w:[ 10 12 -1 9 ]
  _GGAND4x8 #(10) g15 (.I0(x4), .I1({8{w36}}), .I2({8{w37}}), .I3({8{s2}}), .Z(w39));   //: @(407,247) /sn:0 /w:[ 1 1 1 5 0 ]
  //: IN g20 (s2) @(269,488) /sn:0 /w:[ 29 ]
  //: joint g31 (s0) @(204, 124) /w:[ 26 28 -1 25 ]
  //: joint g39 (s0) @(204, 206) /w:[ 18 20 -1 17 ]
  //: joint g43 (s2) @(277, 255) /w:[ 4 6 -1 3 ]
  //: joint g48 (s2) @(277, 345) /w:[ 22 21 -1 24 ]
  //: OUT g17 (y0) @(655,222) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g25 (.I(s1), .Z(w3));   //: @(307,65) /sn:0 /w:[ 23 0 ]
  //: joint g29 (s2) @(277, 144) /w:[ 16 18 -1 15 ]
  _GGNBUF #(2) g42 (.I(s1), .Z(w37));   //: @(309,250) /sn:0 /w:[ 9 0 ]
  //: joint g52 (s1) @(243, 293) /w:[ 4 6 -1 3 ]
  //: IN g5 (x5) @(66,263) /sn:0 /w:[ 0 ]
  _GGAND4x8 #(10) g14 (.I0(x6), .I1({8{w31}}), .I2({8{s1}}), .I3({8{s2}}), .Z(w34));   //: @(407,330) /sn:0 /w:[ 1 1 0 23 0 ]
  //: joint g44 (s0) @(204, 245) /w:[ 14 16 -1 13 ]
  //: joint g47 (s0) @(204, 336) /w:[ 6 8 -1 5 ]
  //: joint g21 (s0) @(204, 372) /w:[ 2 4 -1 1 ]
  _GGNBUF #(2) g24 (.I(s0), .Z(w1));   //: @(306,49) /sn:0 /w:[ 29 0 ]
  //: joint g36 (s2) @(277, 179) /w:[ 12 14 -1 11 ]
  //: joint g23 (s2) @(277, 387) /w:[ 26 25 -1 28 ]
  _GGNBUF #(2) g41 (.I(s0), .Z(w36));   //: @(308,240) /sn:0 /w:[ 15 0 ]
  //: joint g40 (s1) @(243, 211) /w:[ 12 14 -1 11 ]
  //: IN g0 (x0) @(61,78) /sn:0 /w:[ 0 ]
  //: joint g22 (s1) @(243, 381) /w:[ 26 25 -1 28 ]
  _GGNBUF #(2) g26 (.I(s2), .Z(w4));   //: @(307,81) /sn:0 /w:[ 19 0 ]
  _GGNBUF #(2) g35 (.I(s2), .Z(w13));   //: @(313,182) /sn:0 /w:[ 13 0 ]
  //: joint g45 (s1) @(243, 252) /w:[ 8 10 -1 7 ]
  _GGNBUF #(2) g46 (.I(s0), .Z(w31));   //: @(315,327) /sn:0 /w:[ 7 0 ]
  _GGAND4x8 #(10) g12 (.I0(x5), .I1({8{s0}}), .I2({8{w22}}), .I3({8{s2}}), .Z(w24));   //: @(407,290) /sn:0 /w:[ 1 11 1 0 0 ]
  //: IN g18 (s0) @(191,431) /sn:0 /w:[ 0 ]
  //: joint g30 (s1) @(243, 128) /w:[ 20 22 -1 19 ]
  //: joint g33 (s0) @(204, 167) /w:[ 22 24 -1 21 ]
  //: joint g49 (s1) @(243, 337) /w:[ 1 2 -1 24 ]

endmodule
//: /netlistEnd

//: /netlistBegin adder
module adder(res, b0, a0, sign);
//: interface  /sz:(98, 48) /bd:[ Li0>a0[7:0](16/48) Li1>b0[7:0](32/48) Ro0<res[7:0](16/48) Ro1<sign(32/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output sign;    //: /sn:0 {0}(36,333)(36,472)(63,472)(63,453)(80,453){1}
output [7:0] res;    //: /sn:0 {0}(#:609,476)(609,537)(574,537)(574,550)(589,550){1}
input [7:0] a0;    //: /sn:0 {0}(#:133,79)(143,79)(#:143,138){1}
input [7:0] b0;    //: /sn:0 {0}(#:495,91)(504,91)(#:504,116){1}
supply0 w52;    //: /sn:0 {0}(710,160)(710,150)(652,150)(652,230){1}
wire w32;    //: /sn:0 {0}(495,231)(495,159)(158,159)(158,144){1}
wire w45;    //: /sn:0 {0}(440,231)(440,146)(509,146)(509,122){1}
wire w46;    //: /sn:0 {0}(49,233)(49,200)(469,200)(469,122){1}
wire w38;    //: /sn:0 {0}(411,331)(411,411)(604,411)(604,470){1}
wire w51;    //: /sn:0 {0}(684,330)(684,340)(669,340)(669,216)(563,216)(563,231){1}
wire w37;    //: /sn:0 {0}(280,234)(280,178)(138,178)(138,144){1}
wire w34;    //: /sn:0 {0}(595,331)(595,337)(585,337)(585,216)(479,216)(479,231){1}
wire w21;    //: /sn:0 {0}(495,331)(495,439)(594,439)(594,470){1}
wire w43;    //: /sn:0 {0}(697,230)(697,147)(539,147)(539,122){1}
wire w31;    //: /sn:0 {0}(524,231)(524,137)(519,137)(519,122){1}
wire w28;    //: /sn:0 {0}(668,330)(668,429)(574,429)(574,470){1}
wire w23;    //: /sn:0 {0}(194,333)(194,369)(624,369)(624,470){1}
wire w24;    //: /sn:0 {0}(107,334)(107,381)(634,381)(634,470){1}
wire w36;    //: /sn:0 {0}(309,234)(309,162)(499,162)(499,122){1}
wire w41;    //: /sn:0 {0}(107,234)(107,187)(118,187)(118,144){1}
wire w25;    //: /sn:0 {0}(20,333)(20,402)(644,402)(644,470){1}
wire w35;    //: /sn:0 {0}(511,331)(511,341)(496,341)(496,242)(410,242)(410,221)(395,221)(395,231){1}
wire w40;    //: /sn:0 {0}(136,234)(136,192)(479,192)(479,122){1}
wire w30;    //: /sn:0 {0}(210,333)(210,343)(195,343)(195,219)(91,219)(91,234){1}
wire w22;    //: /sn:0 {0}(280,334)(280,391)(614,391)(614,470){1}
wire w44;    //: /sn:0 {0}(608,231)(608,137)(529,137)(529,122){1}
wire w49;    //: /sn:0 {0}(411,231)(411,166)(148,166)(148,144){1}
wire w27;    //: /sn:0 {0}(194,233)(194,184)(128,184)(128,144){1}
wire w33;    //: /sn:0 {0}(579,331)(579,455)(584,455)(584,470){1}
wire w48;    //: /sn:0 {0}(579,231)(579,155)(168,155)(168,144){1}
wire w29;    //: /sn:0 {0}(296,334)(296,344)(281,344)(281,218)(178,218)(178,233){1}
wire w47;    //: /sn:0 {0}(668,230)(668,172)(178,172)(178,144){1}
wire w42;    //: /sn:0 {0}(123,334)(123,344)(108,344)(108,218)(4,218)(4,233){1}
wire w50;    //: /sn:0 {0}(20,233)(20,159)(108,159)(108,144){1}
wire w26;    //: /sn:0 {0}(223,233)(223,150)(489,150)(489,122){1}
wire w39;    //: /sn:0 {0}(427,331)(427,341)(412,341)(412,219)(264,219)(264,234){1}
//: enddecls

  //: OUT g51 (res) @(586,550) /sn:0 /w:[ 1 ]
  adder g50 (.a(w45), .b(w49), .cin(w35), .cout(w39), .s(w38));   //: @(379, 232) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  adder g53 (.a(w43), .b(w47), .cin(w52), .cout(w51), .s(w28));   //: @(636, 231) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  assign res = {w25, w24, w23, w22, w38, w21, w33, w28}; //: CONCAT g39  @(609,475) /sn:0 /R:3 /w:[ 0 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:1
  adder g43 (.a(w31), .b(w32), .cin(w34), .cout(w35), .s(w21));   //: @(463, 232) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  adder g48 (.a(w44), .b(w48), .cin(w51), .cout(w34), .s(w33));   //: @(547, 232) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  assign {w46, w40, w26, w36, w45, w31, w44, w43} = b0; //: CONCAT g42  @(504,117) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: IN g52 (b0) @(493,91) /sn:0 /w:[ 0 ]
  adder g44 (.a(w36), .b(w37), .cin(w39), .cout(w29), .s(w22));   //: @(248, 235) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  //: IN g47 (a0) @(131,79) /sn:0 /w:[ 0 ]
  adder g41 (.a(w26), .b(w27), .cin(w29), .cout(w30), .s(w23));   //: @(162, 234) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  //: OUT g40 (sign) @(77,453) /sn:0 /w:[ 1 ]
  adder g54 (.a(w46), .b(w50), .cin(w42), .cout(sign), .s(w25));   //: @(-12, 234) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  adder g45 (.a(w40), .b(w41), .cin(w30), .cout(w42), .s(w24));   //: @(75, 235) /sz:(64, 98) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>1 Bo0<0 Bo1<0 ]
  assign {w50, w41, w27, w37, w49, w32, w48, w47} = a0; //: CONCAT g46  @(143,139) /sn:0 /R:1 /w:[ 1 1 1 1 1 1 1 1 1 ] /dr:0 /tp:0 /drp:0
  //: GROUND g49 (w52) @(710,166) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

