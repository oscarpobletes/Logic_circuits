//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg a1;    //: /sn:0 {0}(95,178)(177,178)(177,185)(192,185){1}
reg b1;    //: /sn:0 {0}(94,223)(170,223)(170,201)(192,201){1}
reg a0;    //: /sn:0 {0}(98,61)(162,61)(162,99)(193,99){1}
reg b0;    //: /sn:0 {0}(92,111)(171,111)(171,115)(193,115){1}
wire w6;    //: /sn:0 {0}(453,190)(453,215)(387,215)(387,201)(296,201){1}
wire w7;    //: /sn:0 {0}(413,191)(413,204)(402,204)(402,185)(296,185){1}
wire w3;    //: /sn:0 {0}(400,90)(400,99)(297,99){1}
wire w2;    //: /sn:0 {0}(428,93)(428,103)(413,103)(413,115)(297,115){1}
//: enddecls

  //: LED g8 (w7) @(413,184) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g4 (a1) @(78,178) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: comment g13 @(464,176) /sn:0
  //: /line:"One"
  //: /end
  //: SWITCH g3 (b0) @(75,111) /sn:0 /w:[ 0 ] /st:0 /dn:1
  semiadder g2 (.a0(a1), .b0(b1), .C(w7), .s0(w6));   //: @(193, 169) /sz:(102, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  //: SWITCH g1 (a0) @(81,61) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: comment g11 @(444,76) /sn:0
  //: /line:"One"
  //: /line:""
  //: /end
  //: comment g10 @(387,57) /sn:0
  //: /line:"Both"
  //: /end
  //: LED g6 (w3) @(400,83) /sn:0 /w:[ 0 ] /type:0
  //: LED g9 (w6) @(453,183) /sn:0 /w:[ 0 ] /type:0
  //: LED g7 (w2) @(428,86) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g5 (b1) @(77,223) /sn:0 /w:[ 0 ] /st:0 /dn:1
  semiadder g0 (.a0(a0), .b0(b0), .C(w3), .s0(w2));   //: @(194, 83) /sz:(102, 48) /sn:0 /p:[ Li0>1 Li1>1 Ro0<1 Ro1<1 ]
  //: comment g12 @(403,156) /sn:0
  //: /line:"Both"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin semiadder
module semiadder(C, s0, b0, a0);
//: interface  /sz:(102, 48) /bd:[ Li0>b0(32/48) Li1>a0(16/48) Ro0<s0(32/48) Ro1<C(16/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output s0;    //: /sn:0 {0}(340,79)(289,79)(289,102)(274,102){1}
input a0;    //: /sn:0 {0}(79,124)(114,124){1}
//: {2}(118,124)(128,124){3}
//: {4}(132,124)(156,124)(156,167)(191,167){5}
//: {6}(130,122)(130,101)(184,101){7}
//: {8}(116,122)(116,64)(184,64){9}
input b0;    //: /sn:0 {0}(89,175)(118,175){1}
//: {2}(122,175)(126,175)(126,172)(136,172){3}
//: {4}(140,172)(191,172){5}
//: {6}(138,170)(138,106)(184,106){7}
//: {8}(120,173)(120,163)(126,163)(126,69)(184,69){9}
output C;    //: /sn:0 {0}(267,170)(212,170){1}
wire w8;    //: /sn:0 {0}(253,99)(220,99)(220,67)(205,67){1}
wire w5;    //: /sn:0 {0}(253,104)(205,104){1}
//: enddecls

  //: joint g8 (a0) @(116, 124) /w:[ 2 8 1 -1 ]
  _GGAND2 #(6) g4 (.I0(a0), .I1(b0), .Z(C));   //: @(202,170) /sn:0 /w:[ 5 5 1 ]
  //: OUT g3 (C) @(264,170) /sn:0 /w:[ 0 ]
  //: OUT g2 (s0) @(337,79) /sn:0 /w:[ 0 ]
  //: IN g1 (b0) @(87,175) /sn:0 /w:[ 0 ]
  //: joint g11 (b0) @(138, 172) /w:[ 4 6 3 -1 ]
  //: joint g10 (b0) @(120, 175) /w:[ 2 8 1 -1 ]
  _GGAND2 #(6) g6 (.I0(!a0), .I1(b0), .Z(w8));   //: @(195,67) /sn:0 /w:[ 9 9 1 ]
  //: joint g9 (a0) @(130, 124) /w:[ 4 6 3 -1 ]
  _GGOR2 #(6) g7 (.I0(w8), .I1(w5), .Z(s0));   //: @(264,102) /sn:0 /w:[ 0 0 1 ]
  _GGAND2 #(6) g5 (.I0(a0), .I1(!b0), .Z(w5));   //: @(195,104) /sn:0 /w:[ 7 7 1 ]
  //: IN g0 (a0) @(77,124) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

