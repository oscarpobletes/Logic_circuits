//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "LG_prime_numbers.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg x1;    //: /sn:0 {0}(502,467)(410,467)(410,472)(400,472){1}
//: {2}(398,470)(398,440){3}
//: {4}(400,438)(410,438)(410,433)(502,433){5}
//: {6}(398,436)(398,400){7}
//: {8}(400,398)(458,398)(458,397)(509,397){9}
//: {10}(398,396)(398,358){11}
//: {12}(400,356)(455,356)(455,355)(507,355){13}
//: {14}(398,354)(398,288)(364,288){15}
//: {16}(398,474)(398,494){17}
reg x3;    //: /sn:0 {0}(189,289)(207,289)(207,343){1}
//: {2}(209,345)(507,345){3}
//: {4}(207,347)(207,385){5}
//: {6}(209,387)(509,387){7}
//: {8}(207,389)(207,420){9}
//: {10}(209,422)(219,422)(219,423)(502,423){11}
//: {12}(207,424)(207,456){13}
//: {14}(209,458)(219,458)(219,457)(502,457){15}
//: {16}(207,460)(207,493){17}
reg x2;    //: /sn:0 {0}(273,289)(297,289)(297,348){1}
//: {2}(299,350)(507,350){3}
//: {4}(297,352)(297,390){5}
//: {6}(299,392)(509,392){7}
//: {8}(297,394)(297,428){9}
//: {10}(299,430)(309,430)(309,428)(502,428){11}
//: {12}(297,432)(297,463){13}
//: {14}(299,465)(309,465)(309,462)(502,462){15}
//: {16}(297,467)(297,492){17}
wire w6;    //: /sn:0 {0}(613,371)(587,371)(587,409)(549,409)(549,428)(523,428){1}
wire L2;    //: /sn:0 {0}(634,368)(676,368)(676,335){1}
wire w2;    //: /sn:0 {0}(613,366)(568,366)(568,392)(530,392){1}
wire w5;    //: /sn:0 {0}(613,361)(566,361)(566,350)(528,350){1}
wire w9;    //: /sn:0 {0}(613,376)(598,376)(598,448)(555,448)(555,462)(523,462){1}
//: enddecls

  //: SWITCH g4 (x1) @(347,288) /sn:0 /w:[ 15 ] /st:0 /dn:1
  //: joint g8 (x1) @(398, 356) /w:[ 12 14 -1 11 ]
  //: SWITCH g3 (x2) @(256,289) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g13 (x2) @(297, 392) /w:[ 6 5 -1 8 ]
  //: SWITCH g2 (x3) @(172,289) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: comment g1 @(172,91) /sn:0
  //: /line:"F2 Example:"
  //: /line:"N  | x3 x2 x1 |F2(x3,x2,x1)"
  //: /line:"0    0   0  0      0"
  //: /line:"1    0   0  1      0"
  //: /line:"2    0   1  0      1"
  //: /line:"3    0   1  1      1"
  //: /line:"4    1   0  0      0"
  //: /line:"5    1   0  1      1"
  //: /line:"6    1   1  0      0"
  //: /line:"7    1   1  1      1"
  //: /line:""
  //: /end
  _GGAND3 #(8) g11 (.I0(x3), .I1(x2), .I2(x1), .Z(w9));   //: @(513,462) /sn:0 /w:[ 15 15 0 1 ]
  //: joint g16 (x2) @(297, 430) /w:[ 10 9 -1 12 ]
  _GGAND3 #(8) g10 (.I0(x3), .I1(!x2), .I2(x1), .Z(w6));   //: @(513,428) /sn:0 /w:[ 11 11 5 1 ]
  //: joint g19 (x2) @(297, 465) /w:[ 14 13 -1 16 ]
  //: joint g6 (x3) @(207, 345) /w:[ 2 1 -1 4 ]
  //: LED L2 (L2) @(676,328) /w:[ 1 ] /type:0
  //: joint g7 (x2) @(297, 350) /w:[ 2 1 -1 4 ]
  _GGAND3 #(8) g9 (.I0(!x3), .I1(x2), .I2(x1), .Z(w2));   //: @(520,392) /sn:0 /w:[ 7 7 9 1 ]
  //: joint g15 (x3) @(207, 422) /w:[ 10 9 -1 12 ]
  //: joint g20 (x1) @(398, 472) /w:[ 1 2 -1 16 ]
  //: joint g17 (x1) @(398, 438) /w:[ 4 6 -1 3 ]
  _GGAND3 #(8) g5 (.I0(!x3), .I1(x2), .I2(!x1), .Z(w5));   //: @(518,350) /sn:0 /w:[ 3 3 13 1 ]
  //: joint g14 (x1) @(398, 398) /w:[ 8 10 -1 7 ]
  _GGOR4 #(10) g21 (.I0(w5), .I1(w2), .I2(w6), .I3(w9), .Z(L2));   //: @(624,368) /sn:0 /w:[ 0 0 0 0 0 ]
  //: comment g0 @(170,23) /sn:0
  //: /line:"Exercise:"
  //: /line:"Design a circuit that shows only prime numbers given the combination x3,x2,x1"
  //: /line:""
  //: /line:"F2=notx3*x2*notx1 V not*x3*x2*x1 V x3*notx2*x1 V x3*x1*x1..."
  //: /end
  //: joint g12 (x3) @(207, 387) /w:[ 6 5 -1 8 ]
  //: joint g18 (x3) @(207, 458) /w:[ 14 13 -1 16 ]

endmodule
//: /netlistEnd

