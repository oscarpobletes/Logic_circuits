//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "B_greater_than_A.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg x1;    //: /sn:0 {0}(558,414)(428,414)(428,422)(418,422){1}
//: {2}(416,420)(416,394){3}
//: {4}(418,392)(428,392)(428,373)(557,373){5}
//: {6}(416,390)(416,340){7}
//: {8}(418,338)(428,338)(428,330)(558,330){9}
//: {10}(416,336)(416,299){11}
//: {12}(418,297)(424,297)(424,286)(560,286){13}
//: {14}(416,295)(416,249){15}
//: {16}(418,247)(428,247)(428,243)(558,243){17}
//: {18}(416,245)(416,207){19}
//: {20}(418,205)(428,205)(428,197)(556,197){21}
//: {22}(416,203)(416,156){23}
//: {24}(418,154)(428,154)(428,145)(549,145){25}
//: {26}(416,152)(416,111)(401,111){27}
//: {28}(416,424)(416,475){29}
reg x0;    //: /sn:0 {0}(558,419)(514,419)(514,430)(504,430){1}
//: {2}(502,428)(502,387){3}
//: {4}(504,385)(514,385)(514,378)(557,378){5}
//: {6}(502,383)(502,348){7}
//: {8}(504,346)(514,346)(514,335)(558,335){9}
//: {10}(502,344)(502,310){11}
//: {12}(504,308)(514,308)(514,291)(560,291){13}
//: {14}(502,306)(502,250){15}
//: {16}(504,248)(558,248){17}
//: {18}(502,246)(502,217){19}
//: {20}(504,215)(510,215)(510,202)(556,202){21}
//: {22}(502,213)(502,157){23}
//: {24}(504,155)(549,155){25}
//: {26}(502,153)(502,111)(493,111){27}
//: {28}(502,432)(502,482){29}
reg x3;    //: /sn:0 {0}(549,125)(285,125)(285,127)(275,127){1}
//: {2}(273,125)(273,110)(252,110){3}
//: {4}(273,129)(273,185){5}
//: {6}(275,187)(556,187){7}
//: {8}(273,189)(273,231){9}
//: {10}(275,233)(558,233){11}
//: {12}(273,235)(273,280){13}
//: {14}(275,282)(285,282)(285,276)(560,276){15}
//: {16}(273,284)(273,319){17}
//: {18}(275,321)(285,321)(285,320)(558,320){19}
//: {20}(273,323)(273,358){21}
//: {22}(275,360)(285,360)(285,363)(557,363){23}
//: {24}(273,362)(273,402){25}
//: {26}(275,404)(558,404){27}
//: {28}(273,406)(273,481){29}
reg x2;    //: /sn:0 {0}(330,110)(337,110)(337,142){1}
//: {2}(339,144)(349,144)(349,135)(549,135){3}
//: {4}(337,146)(337,197){5}
//: {6}(339,199)(349,199)(349,192)(556,192){7}
//: {8}(337,201)(337,237){9}
//: {10}(339,239)(349,239)(349,238)(558,238){11}
//: {12}(337,241)(337,283){13}
//: {14}(339,285)(349,285)(349,281)(560,281){15}
//: {16}(337,287)(337,334){17}
//: {18}(339,336)(349,336)(349,325)(558,325){19}
//: {20}(337,338)(337,375){21}
//: {22}(339,377)(345,377)(345,368)(557,368){23}
//: {24}(337,379)(337,406){25}
//: {26}(339,408)(349,408)(349,409)(558,409){27}
//: {28}(337,410)(337,486){29}
wire w6;    //: /sn:0 {0}(579,240)(594,240){1}
wire [3:0] w4;    //: /sn:0 {0}(#:555,140)(638,140){1}
//: {2}(642,140)(722,140)(#:722,121){3}
//: {4}(640,138)(640,119){5}
wire w23;    //: /sn:0 {0}(765,281)(765,306)(703,306){1}
wire w22;    //: /sn:0 {0}(631,241)(631,299)(682,299){1}
wire w12;    //: /sn:0 {0}(682,309)(594,309)(594,327)(579,327){1}
wire w2;    //: /sn:0 {0}(577,194)(667,194)(667,294)(682,294){1}
wire w29;    //: /sn:0 {0}(682,319)(642,319)(642,411)(579,411){1}
wire w9;    //: /sn:0 {0}(682,304)(596,304)(596,283)(581,283){1}
wire w26;    //: /sn:0 {0}(682,314)(619,314)(619,370)(578,370){1}
//: enddecls

  //: joint g8 (w4) @(640, 140) /w:[ 2 4 1 -1 ]
  //: SWITCH g4 (x0) @(476,111) /sn:0 /w:[ 27 ] /st:0 /dn:1
  //: joint g37 (x2) @(337, 377) /w:[ 22 21 -1 24 ]
  //: joint g34 (x1) @(416, 338) /w:[ 8 10 -1 7 ]
  _GGAND4 #(10) g13 (.I0(!x3), .I1(x2), .I2(!x1), .I3(!x0), .Z(w2));   //: @(567,194) /sn:0 /w:[ 7 7 21 21 0 ]
  //: SWITCH g3 (x1) @(384,111) /sn:0 /w:[ 27 ] /st:0 /dn:1
  //: SWITCH g2 (x2) @(313,110) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g1 (x3) @(235,110) /sn:0 /w:[ 3 ] /st:0 /dn:1
  _GGAND4 #(10) g16 (.I0(x3), .I1(x2), .I2(!x1), .I3(!x0), .Z(w12));   //: @(569,327) /sn:0 /w:[ 19 19 9 9 1 ]
  //: joint g11 (x1) @(416, 154) /w:[ 24 26 -1 23 ]
  //: joint g28 (x3) @(273, 282) /w:[ 14 13 -1 16 ]
  //: joint g10 (x2) @(337, 144) /w:[ 2 1 -1 4 ]
  //: joint g32 (x3) @(273, 321) /w:[ 18 17 -1 20 ]
  //: joint g27 (x0) @(502, 248) /w:[ 16 18 -1 15 ]
  _GGAND4 #(10) g19 (.I0(x3), .I1(x2), .I2(x1), .I3(!x0), .Z(w29));   //: @(569,411) /sn:0 /w:[ 27 27 0 0 1 ]
  //: joint g38 (x0) @(502, 385) /w:[ 4 6 -1 3 ]
  //: LED g6 (w4) @(722,114) /sn:0 /w:[ 3 ] /type:3
  //: joint g9 (x3) @(273, 127) /w:[ 1 2 -1 4 ]
  assign w4 = {x3, x2, x1, x0}; //: CONCAT g7  @(554,140) /sn:0 /w:[ 0 0 3 25 25 ] /dr:0 /tp:0 /drp:1
  //: joint g31 (x0) @(502, 308) /w:[ 12 14 -1 11 ]
  //: joint g20 (x3) @(273, 187) /w:[ 6 5 -1 8 ]
  _GGAND4 #(10) g15 (.I0(x3), .I1(!x2), .I2(!x1), .I3(x0), .Z(w9));   //: @(571,283) /sn:0 /w:[ 15 15 13 13 1 ]
  //: joint g39 (x1) @(416, 392) /w:[ 4 6 -1 3 ]
  //: joint g43 (x1) @(416, 422) /w:[ 1 2 -1 28 ]
  //: joint g29 (x2) @(337, 285) /w:[ 14 13 -1 16 ]
  //: joint g25 (x2) @(337, 239) /w:[ 10 9 -1 12 ]
  _GGOR6 #(14) g17 (.I0(w2), .I1(w22), .I2(w9), .I3(w12), .I4(w26), .I5(w29), .Z(w23));   //: @(693,306) /sn:0 /w:[ 1 1 0 0 0 0 1 ]
  //: joint g42 (x0) @(502, 430) /w:[ 1 2 -1 28 ]
  _GGAND4 #(10) g14 (.I0(x3), .I1(!x2), .I2(!x1), .I3(!x0), .Z(w6));   //: @(569,240) /sn:0 /w:[ 11 11 17 17 0 ]
  //: LED g5 (w4) @(640,112) /sn:0 /w:[ 5 ] /type:1
  //: comment g44 @(254,510) /sn:0
  //: /line:"We could factor or reduce with disjunctive normal form"
  //: /end
  //: joint g36 (x3) @(273, 360) /w:[ 22 21 -1 24 ]
  //: joint g24 (x3) @(273, 233) /w:[ 10 9 -1 12 ]
  //: joint g21 (x2) @(337, 199) /w:[ 6 5 -1 8 ]
  //: joint g41 (x3) @(273, 404) /w:[ 26 25 -1 28 ]
  //: joint g23 (x0) @(502, 215) /w:[ 20 22 -1 19 ]
  //: joint g40 (x2) @(337, 408) /w:[ 26 25 -1 28 ]
  //: comment g46 @(636,159) /sn:0
  //: /line:"4 bits"
  //: /end
  //: comment g45 @(258,530) /sn:0
  //: /line:"Or optimize with Karnaugh maps"
  //: /end
  //: joint g35 (x0) @(502, 346) /w:[ 8 10 -1 7 ]
  //: joint g26 (x1) @(416, 247) /w:[ 16 18 -1 15 ]
  //: joint g22 (x1) @(416, 205) /w:[ 20 22 -1 19 ]
  //: comment g0 @(26,11) /sn:0
  //: /line:"Determine if B>A given the next table:"
  //: /line:""
  //: /line:"B= b1 b0"
  //: /line:"A= a1 a0"
  //: /line:""
  //: /line:"      b1  b0  a1  a0"
  //: /line:"N |  x3  x2  x1  x0 | B>A"
  //: /line:"0    0   0   0    0    0"
  //: /line:"1    0   0   0    1    0"
  //: /line:"2    0   0   1    0    0"
  //: /line:"3    0   0   1    1    0"
  //: /line:"4    0   1   0    0    1"
  //: /line:"5    0   0   1    1    0"
  //: /line:"6    0   1   0    1    0"
  //: /line:"7    0   1   1    1    0"
  //: /line:"8    1   0   0    0    1"
  //: /line:"9    1   0   0    1    1"
  //: /line:"10   1   0   1    0    0"
  //: /line:"11   1   0   1    1    0"
  //: /line:"12   1   1   0    0    1"
  //: /line:"13   1   1   0    1    1"
  //: /line:"14   1   1   1    0    1"
  //: /line:"15   1   1   1    1    0"
  //: /end
  _GGAND4 #(10) g18 (.I0(x3), .I1(x2), .I2(!x1), .I3(x0), .Z(w26));   //: @(568,370) /sn:0 /w:[ 23 23 5 5 1 ]
  //: joint g12 (x0) @(502, 155) /w:[ 24 26 -1 23 ]
  //: joint g33 (x2) @(337, 336) /w:[ 18 17 -1 20 ]
  //: joint g30 (x1) @(416, 297) /w:[ 12 14 -1 11 ]
  //: LED Y (w23) @(765,274) /w:[ 0 ] /type:0

endmodule
//: /netlistEnd

